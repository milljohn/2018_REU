// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0.1
// ALTERA_TIMESTAMP:Thu Jun  4 11:11:14 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BDAyGi+G2g/enYIqSbzDYy0k+lopOqVHOeWgidqDys/8b7wGAtR9HAStcOIaNJeW
O+tCm+TAlsQuK/4xNBUVylDt89jLIOokBGBz/2Yfe4zblG+HR1u6/7XWur8j1BJt
JcXS2WF7mWhglROLepK4W8K7WcmECyBrQw9tBH0jpv0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20672)
8GlmdBoEfKNMvAzL2uIxBsltZjdaOmfJGeOUCPSHe1Pudopzeyeiv8nfivxpFvMG
jdYvhTAEEqbMoKpiDRL+fO5nToRdkHWHSDYPltCYS8pFzZGcbnVCPQtB6GqrD3y3
ewjnn57+hbgjuGuhJa6KFnTNib/AodmET8NirNn/Z5dvcp94sNmpmgeZr8lCnTcN
nEQo592uYBGkYK+LL7b6WnhRps8kOIIUTqtFOl+KcXOyKyU3h3G34IIhqdWEeGFo
aH8LtIT86H+PEmlo8l+SB93NC5yJZ913p4in+74IChuLoVlQMj4GRLXcbl8Bmhze
qB6pYWiQZfziTdxQeHEabjlKxfj6Dh11Km5xEvmW8S3Mp6NZ4AutXrj8rUWWVuSo
nCso4vVl39VyQSIzzZYYDgDVRxVEMd4ClVE5Y9I5CF1MN4Q44OQ5/+ddXJB12Ztf
eMG24snT3Q263L1B1swfWjcAe7kEnXtZRZePMu2ddfTpp5mzsIapIF9NfrJjZjSM
3hgXxsmXOxhqeHc3hN8+MpY8lw2DTpRpXRKMGpi9j+XGgg8el4ZsGRZQra5a5Y5g
t/0XF0gE9SUuGFnN462+pl71k3naiLpF5ItY/pxT0YH9T3Pzj8lMahxL0gg5j9rM
k2iYjWruzBARyACqjloNjA8DgjAIb5U/BMrzrQ3RA+PDqK0fDnmzPLGzvGhsF0un
LrwhT6Rca8IilEb0iouE4CEPLRRVjxKkBzx9uPAED1aODL3OzITUAs5tuhfqslpP
vI+UsUKtiX/GmmK+EkDTtp4ubAZjor6BA65cjdq42IJ4ktwf2MuRuHF5EOMC2Zdo
I21+3XqfnRme6840KM/95pUhpFF6k5otJuK7p1PWa3j0ETTumFYck7UcsEkqjTd2
oShzvcbGikIym2gp9cnfmu/p7c4LjITVYq5TvDHzamKMDxg6zx6C8kxbTUG43Jvm
y2qwzSU+0jd6l7LPy+jYpwnDmS0Bvk7cjQ8Vg9zwHBx40WIQ76aQ5FgksGSDPpA9
VOukqDgzitL9K2yuW2uH6exsmE4qK78q6m7Wj2F3AcJSkAmbo+hkzmN/EfozJwGJ
YtdXaStQz/ISoPUzLgMOlFqNmwBm0O3gyfnCkK1Aw1FLovhDyJJMUqxzffKEcuVX
BKBXqFJUsV7MxS29CryOxYBvAq73VoZAYp3bYwFu6B3cEUcsIEoxYZsKium3fusi
ILMc820pfG+C9/AGQigj+kMvYJdffqKYsKM4jd2KNhSTZSJiKLRy5Fijcv+PBkK7
oSrwRVjaZKPlt9d1N3GOZ3cA29Ks50i2UY3S/W+OzBfnGldcoiyoR+6EiUymMb4M
FnJrDS03iiCPdsZ56kEgQnf4Jaqiv6pm4yuCe87OQAewmeaVfMflSsbbbKfyzFTr
gquv0q+P5OS8lvetSA+iQp41sR6UlUuoKF8GCKC9sKIw+DZmVFzSOOGtavwF2xBE
JbZEvQx5AgIZ6Or/Yj9SUFgwRkJp907yeYKLmAqObbGKDDrzf1kRzGJRSoJHirxK
f0t+HMxre/YU1L3DhPTduD07TgDlHdZ67a2f+g7ip1GNDqCW+OiEdNN38yoN/IV8
OCBgXwmnwV6dDYM/gd2s00Dvh5dB/shlVrwHfgwCHJ2fwXsEp6oq5UT//+mnZznU
xB6PMtJKN+un6O8O21dXx8J4g4ceWtgTXf1QbKhMaWPY+ypEbe7JjNfVhQEiTGIn
6DSpOCZfqoTXdz7MdjHCrKhn7xKP/XoggBtHcbM447tmp2RQRKTtpTg5WofGPsj8
iDLcl/J14zOA5QjTlMQ5vMdPXyyNYMdYN1AwWip0zVnNqggqSTtbGpM8WPDduOo7
WIRRJkerpHhRO7sD2TYqN1mg/MOABpOUna+H4KMMwHFldFZ/EzwWgXnzfY/G+Qb4
KEBdvf6cW2mw4bLLd4Xh6wJ715lxy7wF4gtndn9QjWNkpAtHMiphqetV2UqxuhB8
xqBzesupNrxOjvy8vvPCi6tZFMkOaUWiziKLfkhNYbfzeeS/hQyV/Jk0R+zxN50M
dHg3FOxSBLUhNa0r4e77IS1CJ58hc94wiKnVRWqQq8x7xwbj+DwY9uL9sNa/e0fj
1T1GTR4RSr6Kb8zPekGzoNvvhWQ2gHwWbdEJhDvYsyvfGGe4e7UsB3VG7+GF2FYD
2UoX3yFChH0JSXOGN3hvR3l8PtyEsRfCBUwHPA/vzv3yM8gBw84cajdeG/SCDO7m
QPohMuY6xvNy9HBMzjjucGoaFMVcwZEMZ18FxuuugZrtJjwbrN/ZgLMcfpeneYn7
c7HB/RmDtPSj2d4KSmXGmP/NgO+fJb4k0L9Rgy7Ie5xSWrz8qjXW+urOpjHts8XI
vAdklYktTX71jzNczcBnJyvleWdngllOJ1S6SMeT4O42HEiweZh13wXJ+DTpjcCX
ryt/gzRQ6nby3lGjI6YM86Qiy+nxnl6d7ImPLYwDvq/MwjTnCVRaOWiu4ftPdLEG
pC7Qmz0Rl8FggJLSX65hQfHc72OUbGeHpGP5QdM+phMRdvfhXDjOU1zbGrftHCLB
9K14dqdbK6I6KrQF0JZajMnCC+WcCAQuWMp3nPW4mX3Ir9jQGPPbt3nkHlgscQoX
k43aXmVP//VvME6BNixfbMr4TV+cAIrGvNPZ8RESqccSJXybTv+VUUk14OTu1qzg
YRuE10DXLGszDpdqDp/2XqAMYglH1dwk7IB0rruOiFM6tgkIeGwqnmMU1dZnxuhP
q0PQ7WJg9ikkUeR2JRf0ulwZTgL2QGDQhQP9RhGy4toH+9ULQ9mtiE+5QMlwFexZ
bcsYfquHlEBoaBXXlHNdYMd7v3wrL6u+7qC71oTNIQacfpBPzD5IIQis7y/ArnpX
x1vo/N5ACPrCBSrNr4QsVmQzfaa3q9wsgs10a60MmFeKxqIWZAjx0ToM7eOMoGj4
xcX2ZE2fRIwe+cnqjJfc9b29sb+9mBeu/l3TGNojqRmb7cInmJzXYK6JDx0b5LuP
cDYUFa5WXf25Aa22uwD4vbVqz5wjsBqURKNUWDUk6/DanzGpO5vHKD/ZhGF7PI3K
9eYi4bHYAO21Aq3WXsFLVHEE3ujKMLwC6A/T8xC/SzTwvKU8bWnSJkHraBQvNTuz
iceBQKJsJfWjMuLVtzeYLb6lfkUVGxhorjI5PgB2wBuHBJOfMH3hjI0JUP12i+8/
HktW53BKt8Fw4etYjLwH1u1UGZaIskiX471kTsuyNveM4xL62RMBUPMJeENAhi/V
XFll740a0znHQ3j1nMYSWmIcsiHtbvM4/qaZX+ctgJcKo7cztEt3Rs3lgygqVej/
PPvoaE53VAZWQFpDbuHVOUrelASFwvRqKjlNr0uhE9ErcO0YA1KSEY1f76fIHoJI
yAURJr1qxiwLj3si9K53wlYxmrplWG2K6h0G62Fy1Hhzjt/Jc1ePNT3SdCU669rR
hP+yk8ZSKoBXXGwcvvQahf5Df/8p8aq/Pkf780KGH0Rhb6dVxq/R0lQvrLQpo+nu
+Pk+xWKB0jAN4HgF8HIjjwkdaend3Cv/mAneqEq/UuEtmZdg4Pbe9LBF/GySr9Mg
R91Gvgey5PhwaWuRMCaeZUeMMnsBjp2VYQHFk6K2QxN79VR4QFgsS5X2n30ysU7b
S0yEeIsUWsSFygWuWdqcNWHLSxzlm1gldnzG3KfJY/TEbzbUQMDHz0pK9rkPCjNN
/2FoOYgr2JR+lNQitQvZIu1GkWG7qzBhvgDLOTAT11ArT6Wc2xXqjf/GkSx92j8y
JCg1xTMyFS9vl6TbI/w06+cL6xiPwUXtotpC2SvBEX9z29/SastjqwQf25qsVKhR
VhIdHQVfxi0XQr//MGS41alvP6jm76cyW09XVBW2Ns+oVuJLhWoXc8ABjSCZZG7/
H2MhxZaOrqFsH8IBdvJz34k+QuMiE1ngcBwl6TOyNqsiY5BBMxf6/sSgBRYjU3+2
Z/Hz2295mr5KP6zTmBeG/L5EaHLibwZHjJbNoiUXFFS708BIVkG788vbryh8HV43
jaz6creN2oKbPnKHg+pxSIOx0rmCbyGr5ra0+XbspJH/IbabQ1I6ZY9zEqnpliN7
8HTcyKNsFW/HDPkSNiAP8sg1VmAyW56zsttE4JklU9jLrTP0/NnqQ6hboFIetjBV
zlhkCl1d2SJwrd5O03P1Ptwbq0PDNCRpGaZR9WH7Nac4xPnfwT4XiBLA32jun3Io
l6Bu+WkNgXhpwvsroeETl3p4334hpmZt8ZUkjI1vkHKsRN1GKRN6PGl+3jqFL+vr
9aWy/Wt0w1VLF0LbBlba43tcknW/ZnNfPEBvtXSNoh6ZWPPq7q8P9yEN8/mLoL5D
GX9pK3MnW0jR8iPiRLiILd+UrRXzBXjMLmN6Hqd1VSsAJvH4tRtXHVW1GVALYwfm
9avmiSyUGJJibqHmatpUu8IfmZQpP/k6L3MNUtCK2xf/AyWJgClzgd2o+iv71fzJ
Y/LCNZ6pK1S5O5nAF51MOdrTzxbtOB8EJ05M/JmTvidW/N0B8tSr9GBHfYINAU8L
fHZO1L+wlTOIgX2aIYUNZAjOmAdO2XvoqeuhaNodHqEZ4ZxU8UWwbiqJwDe6hEKv
xjhEvcDDrlBvFNcU06WaR2oq5RMjcAwQJQ2cKLB60EEko4tZYT+7iPWo22K4HgI6
IwOCpKTSyyJz5ITMFfqT2m5S1uFjMPE7WFpUT3zpeJYqcS/DM3TqAg+TOjmibav/
YFZuLJN7CwO+Z8WjSi+QJ5DVB1Q6CQxg+eIV7EqixvZ0IKVkHyUVk+ydgvvpYNb3
YW7pN9eyBroSyoQ7yrXIQbGFRHlKwUyaRwPYSPDX36wMbqYWm43PUaah3VYlZqHZ
F7V9yb8wxFrAgl1orTpsT2Xuj3sSFFC2tRPwEatdsCRyViWep2CnqxVsFX9mPcnt
P7txQVoa/zk3ZI7blIFDpC0S0QuPBfhwdGKBuhyp6nNTzsYPgvs7jsyhm/rvcRRQ
v+VQaV01gpnW3Yx6oaX4Una2yr9ZEphsWvzev1ExYdmECmOfyY6npP5dY2tQHcau
oAD6GFGhlFscMVd+HGUX4Vbn9BpVjq006PUKDlSiqTm1vbetiWJeGeWCOwv+4NC6
BG+CklnunqEJ8T4nNXwnRdh70B0Oh2Fz1hLL0MpBQZj/mExnPjANpFBLSNTPYuB5
IaZBJIeNdUGo/8ABzMO/sRMmXWJDjI49SMWLJwb1VPYoyKcFSzpI/FEOqK8/L2gI
YvE8mzj5GTbG0r6jGphhOa1jLPSwRPsIgWlX3sVtjgkXirWoM2H6oB41qwkW8tw5
NlGcFj73BAcQ77wxbi2kNnUukaJn+yBJDjoOtKbaKFZJA/7UsPdpNbSleYLw3VKa
uuVpijpTGb+1kfjuayXS+z3fjk/QNxRIdkKX6PyHXVjUFPGgngKamofvVttBfqxl
bE00e5Ha8/PhXVX4t0VXbu7cC82/6PFkQuPRQxizVxz5cC/j8h9I5u8hmDek/9dn
FS6WZmC4CZ8zEpy2xWLwqAEj0q91SSR1djoFMty0ErnPRop16vSiJURnLoIEBAvZ
sWhrDsa04CBOtNs++P4r8EdIFAF70Ej0It2kNkCQ1lq4tAbDicomse+Taf/KHJ9P
kAkZwxm2MQc1Pfh0HclNQUHVj9/pO0rJlqWYA8584abDZJRAxj5cMoCQNR5kS4y0
GFbfpS53ui1A/2lKY9Gr3c60IDCwh3sepTIAZchniQRt8A+LifILcrChic5tOzv5
xSql3DBKu2gWBzqBg0Y3LLRzLkszW7+CHAdE7zYE4NM7ooitFx7/lWTD8I8sDxpa
H2S544CLNJwPc7tR58W3oIcSlnS+rrBrWHIwWCMcgUB49fctlzdbzmCcFUyMpUG1
toLvwLapOWI4iyYnMGK2EWd9+xoXPYFu42uxPbF4PLN7te4l4C3jCZp+RtOZ2c+R
PbCIlO5sDofSdOEA3Ub7N7bueHX/7vAOin7IvxFkyfMqwjXkhA/3EkqnzpZvsvGw
OvGdIL2ykf6iSUEjS7zHF9XySSj7H1pOwH33MM3AQUuLNX970gBiN1O6fTL8mjhh
0GId7CHyzEPUf1RPD2v9ZnAvXU7NAY2xmRDRiXa1MTi7aXMLzjb0nVDewYYyjiUj
aWSS+UIcRKz7Mz0C05a++PhBCY8KriNxhTh9eeIZf1EOL+x1PpmyIeZhE1fecrwz
sIo9m0+ynnSkE+PoJ7TiUbhz8xuKu6MiTrrzHKkQRAQPlT2Ugybgs5mKV3RELQ2q
6tpPQVp0u4gqk9OAaIicL5c2IAWoT0LA4nbqALv/mIc+wjb6BUwmSAHHz3NKAPL2
PkteYA4mBBFqZRb3tMvwz+irp49lCMlyA20FZDOeIrxoagFOl0GRcgNrPonr8+Bl
Iz2LNNHcBZNGcXVdwQrGO3uO/zWE3xLqbCGG6BACruDxEGVHB29hfSmBh/FSaxDd
GO22dCRZtdgCwBRZ810Z9dMMklFy5ERhLztQlKj8C2tOTTWLB+9p9xsTtmSEHyTL
ZVOor195L6O7Qur+AJxUHnq+C0NuvAa0EVKxKts9HHEOzd99HKdHWZLCMF0Am5yq
e/6HixsuvoDGrp8/iJnBR9nT/SGjXRftKFSni1bL2qbSZB21mBWh2Wc3sKVoLIz1
xKd5UscE+Y21iypPgzd9h4k5zarG8A9m/uvJ89eaeyPi8R0iN2Dq7Nz46vjtFYn2
VggoFb/YDo5AALrvjk5iH7VJjUegFbnfPPlt6oN0GVuw0Vt563BGdNlK9ehyfUnG
NtpLHV6AuMAhTU+fyoc/YrZfuupGwo18Nu/rqhATvjd1i0zNCl0w6hm5onaLjeR1
mupMZ/MyKuHB7uXbkpHydy1OkSmkxScbOIpuVzBE1b0o0dIruA1folQ5vf5fkM5I
1NOmbzl9q8aIF6Q7ryF0RmjtL6iI+xbJgvj8bIzEYauQiiVgOyZDb26O6eyAjMEC
Ij3jaVx8WUtvND6foZ//g4vARD7qCFTW8voe4orQdEnlbJ2U///TiBsTTCV1BDCz
XhtwcQ9QyJqKus9BpbNjrXyJxnsgVci9QI2fFwvc8KToUKBwWg5SE7vzq7JKxM5d
ijaEVHBAwwNC8r4qUbc+imZqiTPC5VN71GPadCA5XfiT+S93v8W3/bp8WzNgXreJ
pW6vScqFhgq5v9wX/ClN3AO9A2mq2XB4tyzbqSAiQxiRHiK6GH9uICpE4fL1jZKS
elhA9sBCQ3oQ0OoFx13UJcoHzND5DBYdsmhEFuehX1lYte3428TTSdqNdEY/Zc5n
KGSpXjEkEI1lNBII8t5QEpJkAt4ic+cU/elpbNcOi5TxrlH5J3feAHdGsxKiNsxr
D6g4w8dat8SZ5x7nTUWfySXUHjUDogVU3cg2uOCpDDPQ31onfTICtS9u9yLDJGco
9ZK3s6yNl1sjyqt4QKIjG8oJluYIg2iXujKPyC1XJl+GxihTf99LwqBUu5BsJrVQ
qZii+D3p71fIPq2BIRgVe2fiB1H1B2h6bwi/XnUH6759JzjnV6BT9DSDim2VvymT
3FZfuPg7sNRdq0QJYRXQEJch8Z2/+t0T4uZVZGHPdKXz/I0QW2sELfBOKuz9FpYR
fOVBspxQw+jxUIJpX0+eOePds+Rgg14gatYDQDFFzm3QnkS0R80Xa14VlMzxISJr
ydjdK7d+v1+3uSgSrpJMXFHNnXVf9w9Sfi8RkjD49KWpCRD9qsqRKnvmgoWiVnuP
3I09Ed/mgRyVGHF7vpCr6/HEQgncG6179BucYC8OW6R67ArAyBhF32nVbJAn4rAk
gbCt1/xwbcGfc80KiEwcIUQ9Yuu9jfBFk6veP5MwJDIN5kHBoej/ac2uXY9/RsCi
cb3EdgRQCX0kstJZ2pcgUEJJ2TzQefbwXtyHsFKrTifMo4Dm21Nv02+lCCbebsl9
SeoWbmewE/gTT2ixA+WzNewRXFZGwh8Kbf/aR4B7GScNu/3aH/K4zDtKd+vxWmoG
aZcrvV0B1yusKXE+yNxNdNGmZ4pd3pHbjTqQNhnPp0G5jTblYYDKP15ITnTuKQiT
zgGqk/bLWZdLKCkWxT/uEWlIkeHVRUAUIYyL5tBP0090d/oc90M/Pc6OH8OF0Gnu
BXMer67gtPJ4EwW+rab09fILJGL+VRrMMTmdSOGku513avHnOrO9vw6B1WUlBiTg
EKfs7B+SCSsK9Ri8dNFL3iYy4u3vMcpgLGj5ftyVWELiOy9KKJFBDi4Z4PWBuArY
3g4Ya0fIb+MRPIRG90lgaSsVuCQTKjpqbnlDdOzTmOJD0NP+HgQ9QjGu2XEVOH07
I/LC0LlXGnMsc+ZNr6OSQNPZcgGZb+Wo6CgY1JVlDrbPKCZHYx1ctfA+YZjJFHzS
U3BwN5EdBZ2xH2pm3wyHCrKii/z9w+rqPtE2Ebwu5s86gOrbA8nE5oVQOyFzeSOM
0pf1mHU6F+DetqqiDvratawgMBCXUn96hziHFR0t7dx2f+CMo1q+cBP1CK069qxF
OaXtAWbZlo4nRRc61e1Gcc5Yey87HdOOe8KFnufZ/HkU2MY5YPiTXZ3118Td3F0U
X5H6MIVxj9JIaa/oBYsBQ1S3Qybp+DU4FEzAsuMWJu5I1WLhiXeKB0Zd05MqlQJO
dAENaM8TDr00gh9jszkQ9G5x9bQjOQgBsSWB7C/IBqlHOJzpYMl9ZmWdQOB3+6ef
TOqwAJlniIkDc6q9vjqc/4TWqnEOxbjim8yimgHh+wrwWwOf+J9ryvOBdKAmlwDE
KZxdagxW4/0swx56v8p2ShBUTYtyQB3lezgAOqt86wkuiffF8eIGOboAOiEMffuI
tpYbvRHSVaHxDUg6GPiPMA9YMjt2rM3FcOtfjBz5Xu25I5PcZark8LCx/dDOncIW
/gEWZuxv8WVYCqi7OHNYSaS4xhKlaaMcgaPh2hSFwnjTBYRvLd1EmgqC+31pDLVm
6ly6E34RSct+1Bmw0BiywegisqgI/2JM5d3s2IEITIpjEJDAIhyv9tjaqlYx5B7+
K2RPRTm7efZDT9mj3iXklY1+pbq9wh1b/82JmO3CqCoU/Ij6BU2RStyhU8YQQmGL
5RtZgx+O+FiigQZwT4OI0gXETn2Lms61da3vvVXnYltKLicWgKJuJBa1fvdYITc9
1YH52yoMA21NuWsPTV8fRWvgJzCofep5bKc1te5Bkcx5bZ3Slc5TUIm7YZRqVZLm
Hmve0BQd6Da5duay/jdwy206tYla46JrnN+X8UxgjKMdauIi8hR7MXQ1dOvGwl8t
fnB9NK+xT+Kwx1QYL5EXkQe+T+A+LMhwBoCy8Tvlm97Wiq5db3xvRlv+ac1jadWz
mmih5wmPpDhqKJPe3x8b+FLjqefQh471gh6V79UQJ5PWIoonnp6inm2qhb+Cketn
j01WO4wZm2HObjpJpJD/IOlO4Zlh1zODa6WyhsHCieqJismkzxsAOf0SVebDyCKf
m4k9QHpaIscz74q62vHOCMFZI9zLiV4lIR5wnzBo5OayCS+/kK+mVW/MyW5iWppo
28wvQkOO/gopX8qWI95CWK4hs/o7p86XI/QeG9soGWqrn3fGln5eNLWt48hRN1eE
S1ofXvIEWV773X/53XlVHmX6xwKROy/J8sk+1jTyf32r+awKw72Tjd5tVhRhHmeL
wunQ/sY64TX6vnI7Sd4bsoUolz+7R9jCTBylEOvFcXiXw/P+Hvy/PMo4MQpB99w9
TxRvF8mBOljRaZ/vN7YuEfMlZx2S1u8IrDeqngH90K0369ycIEinrw5tHE26kVoX
uN1Ld+cdi5syTi37swrbvdgMB74ooL8jckMz2XyLG5U+ab0/s79/KNFNTNt6I0yK
o6aQ95B9QypS1E4aZt5JdjuxAnwiqi4VgNY0EtthRkwMi9DcN3L8aaAumkf21ZaA
vgLRjAeSifVCmP25S6qVFZrr9HU+qW1LeQ11D3odrbdXaAHtK67Sky7CXIB3NwZF
bOsL7wil3YydnejYopX55IzajdvEK1DvK6VgZJI7WncaFpyEsEtc6cfwat9xDjCf
9mEAnlORBFYdgpiXHI40dsJk430Q/WWNbrFU03jZZ4mbfJJD/natKfv8sooLMukS
579+xliU3JDmEeRraDVRVkZyoKqaYMKps5ZRKawpyDn/c3BMbylyklrHxGH8N+PQ
RKkGZ2vCcxfFbdOwmghTwKrL1cu5Dc6ekjxRcinieOdpwF2lBJdzXQ9c2k051Iwn
SDqbFmyyd+C0IqePPtY9R1Pw1ixCNVBXWkGVG2X165Mjv0V1MEi/7vA7mwGfdvZZ
TFmYE42CQcE5QkIGg0ayevA22R4kzZ2IXE+pnD+fqaKaehFj31pGsqT2kvKJ5dn2
c4GoGlqWFQcCkq2qyNLMkrzkBahrAmOoeAnmAb8OXt3zlXYKAuGq8kr5NwJmvHSU
vjcBYpM1F4eNnrzlQEhWAVpOI1zPkZJLQBPUtp9RVgCgXSu2OBAJkgb3dXn2xRrC
pIc4PLtT4aumNv5BZsPPuRkJf+xvHkCXnrbci7lWACay1btAxaYwCtbQh3LT4SsB
IdshTDmakLs0PEM+h+ZF7YylWgy4kovFueqLjvF6Uq6zEERvHpzs/xKvvAsAIE3p
24AXWzCLimqKpJmp4sy43dQVCKRLxazdu3al7krmdJ00KpEoJ03aIrJvjHBnm6Er
u/OSYkvLTI85pj8B3ZBPvPBxSnCD+9kUYY1c6pEgss7hq4twPOo2CL6ETKXEyBBO
fwEw+JlpGginwl9M+PfN+vpo9AjbP1eVBFBKXb3qtTx2lwB+4TwpODx+lmlFHieN
x0j/aR5GIM9OUOLI/LL7asVU44HxEB4Ap1uL25m0EZCVpnDnSkf14qDECAEshzoA
ZMyv2itXr+r+cc17mHyfC1hsGRjUKHI7X3WCf8a0XWpeL1Rd6tJaTO1hdyUhyPoF
aMAaPSHc90EabQEcM0lTg6FcUvq2Hi5M5SwnW3Y5Bm0byHH9gsg+ln739/xhGjTB
Wl0ocGBaquPkI4yCFImba3riFw3t7aCkqtR8SIkKYB/k++03kOOApxgHIOh3l/9L
FepmkWzcHGBDd+SUxR4JMAXhjZ/4BmKujE9aXSbFoSnCmvCXmEypUAxD8db6iyfn
xErJ5+fXa5RO0Jnndme9kGpIlnDa0gJWClOtOegRs3g63bWXYJHm8v/uZtxnFUTJ
8A+E3kBUdnTP3KXlEwyT8snh8M/W23X57QnolpPiMsv8A7XbwqHizIQTNn1ETKfC
LyfBG5duw3HJ72rfW8bdQ1jytJc74yJr0xOcHklfNvNrJHCV+rsxslpr3VsLTJCD
Q5p/VRFylOYmJGseofBLk6b1/pDONmwdFqscSSOeTARtXeByQuJ5YUDcUTe+nn8q
hPj7odvc5+ejd8l8GgmoJkW516rupU0mFnbD77M66baL4zsy1aly0qk38JZ4T+bK
PeJFpJczOG9nRuFhae6RC8iY0CDT2bXLJebW6WbeEQhmm0hU9CZVT/h1tIkucLu8
eZ/fj1/qQpFxMaA0FJx1VSpu1/DRjm8jStD9f+BTUzLmAhpTGu/Sv1WGcuhrcmhD
PKl9O+YFVR34/MV2+iVcNkb6U0cruZfD7pMJtASJwGrZimxi/peO3QPepfwpnwkj
85xJXuXm8C49FSJlMQ4vimeGRF3VcDOY+Zvr+gGeP2sqk1LEJthiKGf9xirdcyHX
D2Pa3PSmTpcIwc18ToY2zaiC28QoAexEaV0w4Kjz2lJ2BnttvQlj+/PedYRcDFXc
4LMZDl6li0E77300PmJ+hDf+jFYMS6Pxd4/c9dQvWw9eM0pYbKuNsXQwjmbV+o1g
j+1VvYC4gptn+PzNpxzfm8TjDcrYaY/HdtlmImCtQOUc4xqnXgDaJ8DTAQme21DU
v5Hz5t23Kc+bls8J4J+sf9hQji/ddsRVNQ0enInCrE9SeK1l0FpJlNnvRytKKq2D
52HHzSN2iGvSr38FzBwIGrgsNh/sIfr342bJsDtromEt2GNfu6H1Rdafsc0YB4v1
rQnOR90ZkG8VzJAI7g8ayUjcOXBjhiztG3i9GMCURyp/n8bN4xg9ZkSFnygHMnQl
673mv/iQ7LPCYRtBguY7o0sRZCSfdfdhDWJt9HJUIvSqQ1iwo3rJAajU+BevaLAz
JTMa9idS1Vy5CA95Q6PG0/Q5QnRDg0PL6MIVF/OotGuDxTGo9l4PQyVXuplz4kOl
tGRcb2nz96G3M13L9geVDWQ2IQSr1LTsAyZDZUvgpABnksH8dExvq6vhHeKAvjxB
VUG82vT/BNNhVA2q03Cv7CVZLaz0KdhtYIYgABrIrokVLZK7hPzFsxMx2U0itjNF
yJgbywjkOadlD45NYI0FbxkE6oh5Grsi2QrNiEBmNZJAi8YzcF9igaPD1pXeJdtC
dd8HspuvZTmnCYSoZmd9x3YG6CDs92V6xHYqluXXzmycVtTwTpshDqmM67WZB3BD
CTLuTICTKWUudeTcGKBS9W6USsTyzzJJXwJbGpPDGdcqilUd7UlSKxpjF2xLQ0U8
5ce25WHCckbo6GHxDyA/RWEhLLUb+k+N0yyyaIXXZkNnjqa+x1OwB30/UoJ2tG+d
CDOmYPw9jt7BGLUBhQUWTy1yyiLXRpRi58xkO/W99T2akzQN65JgfS4QEdG2p+NG
L9uAC7OSm92YrDk4mxGgkRqFJYL35RNetGaIbYc2WopC5LT00SM16QVy3yR2kDfv
8xaEAerYsGgS1XZhjK44IYwmuKiydzOywffJ12xuXc0WSSyZoiAXqgpStc8neM+c
0x0EhyhAbHfm6ocQZeOhcs41z9a/w9qPQlf8j7yeFH8WFiATk6H0IzpPuRSuRMaT
bJyFbea7Hjy4Xmoixuiq2t7MLhVsCM0R5hYntSoaTm7SMNY2QiBB62Zch7hNP7kj
l/4z/5ijp2Stp5IqNqFIwTW0N1Afm8AcBjee4lEu76Tg/J7geqJIwkcM4NpZA793
ZpET8WCfgFutgDKEZSPl4v7y0Tna5hPz+ADfaqu6NdXuoCrLqaMYoyQshF0mv8Qv
KoLxQOke3pxwr3MFvmrCT0BhvDefXQvJD+GIKS/nWk6GIRuls0yQvGO/ze9bXNb7
f6VNsptzP9umFZJZUOhAX1S1GJTzKKFag0vLWK2cDA1o5UEWOqRctOQUCsUlYoO3
eEzhPm12rUSJta3U6cg2v6ZPRrkve5XJPM0GEfdfG8+SQEgud8N9kD43PxUiYIer
/tnm39rKlXqzXV2TSSNcueyaxM7t3xIyowB7rqljnSYGJggRMPwieW9dcwLinMwM
Wc86i8pM1KtfAJ/o5mTO5mVcJFLtrPT3RiqGLVv5Btzf3XL1AOz93T6WVBz4EF5N
lDCu3gp5cuGoyYckc6n1+uEbl4B/Shn9rXkanNi5RBSb7ubMEGzvGyz0frfpO75Z
1rha5s6gkGW0/oBegAXxNYsyIcSjJT9WIRrWonJBQgnarzaIR9LmRWh7e7dw2738
VtDLmOIsCCvXyL1mE+Em2uRpgbXICXeo4wQgsTLYIdPqCB/NOmh1cfu77/31SuCN
bWaHvDJusjLnqs2am/raLH8kjuSm95jBr1wTLmRMQlk/VcdhKUGfxmij8Fofsn+J
9ulzZrPYw11eDxg4F1eEpXFJHrQSOs5S3/gcTOF5Rs4TCcZ/ueVcKWgctV/KrlyG
BDK5EC4v427ejvH4hjWw8gD7JWtrisOOL9V7v1QYo7nmAWoeOXMnN8EyrSZnYFPG
2uoSNILXKGnOiGWm8QolQZx9VWhR6y8N1gwaG7vRJFewYzNJG4hE77ZrQfQVx9rb
TMH2o0KO6Gb7U4Gnf6+1De5YEoHGxHCHqubEf/LkQPqT4Bqms/hvYiYcil9+hPdx
HXyCBZfaR7G88SVWTCTDiYWd44mmesFK7ssQ0fv8ySy9j0qlC4uPpwG8UZixqD0G
UnulQTscBDH+orXv65m2FQRXy0MV8/5GXKrSzc3jNfFouItlPqUjU4PIj1w3RzMN
dW2m2bIvW5oDkM6PTJrQUZabH7JryubDqB8F9QKfSip79d4DfRycPI0EAS0zj1c7
6AhAFzkY848P7oAVXtcVH3Zai+5jr3pSwvF3X5ow4vMKKx1bzEXDTSER7ZC3R1KE
/dhhEE4GhDfsU2Igb2YfWv0mS+k3eDPaOvNXQHM75R0XzHPmKr02Obr2Kch/vgoG
hD+GgMkajiWuhysV71AMg4lAeTuA6WRuUO+WR8O/3Z2ene6YTXClMcIE1PhO3BTT
dyWOwyBimh9RKsQGi45legSyVk2uokfzrt0lbmhFLqlmzI1jQapxwzLv4//vgORe
YDQHTTAHe3ust3qNQ7r9+8FmU04AlJCjmlZuBoZ8fkMvQc5h9XjXLVscvZOerBHN
iCVPQVhKA2gJL9X8lkxucGjXhMLnCkzTFfkfHmETNoTm5AWGRew+VJTzU3FUnXED
W/dtnBDvfSrSXPqrGY2fzfSp6U/AjkNRdqibda7pXhrrJ57ANUV5iNFOxeQ40bIi
SP6mzfudt32mPHo4GEiyWJJVxywUa3zTfA/LIqIihN3tM2SG/Eu90KEIXz4NXF3S
G8qPIS+19gQccHRKy1++NGh9LciMvpGwFGo42jtLbdWo60eYAjDg5OdTQkjpgI8A
ABDdrZpT8M+ZiM3QMrSviJSiQ5YReg5D9SQ3Dqd30Ea0Aag5clNGoqKBQ3JG0gpI
n9IQpJgwvSliMipL0wQVyebgesqztfWSNI9zR3GRDZNNkiQ65MlTMQj6sWXXnKZ5
e5VKyFfZepYqDMn3cxdIKXK1v+TBhhulRoi5smpbOq+kOGCb6rgtTp+Eh4TyUA00
iORAXKS10DXn7clrGd7p8swV7BzmFXIX+5MfGrmRKXkjSQcI7alspdbtUeQVwTdA
fyVpxnceyDwbFyVxCEK7fSGzlBJWu6OTzlJ9YI7Nz76e4vPY5UZXWXMS/fpqp0si
2ns+aB6rjqby/oyAX4Evwackr15rm/YO976K6+akK4rFlhj3y28zMeRE0OpBHR84
onaam0mqO93OJDYC2ZcvjzXQRQve0wVs6RwPz8E6Tk9DhQjChjfShPo1LyOdNOju
gULXVtG3AY5dy9FA4zsZaMzKQrXK/4SsnabsNRz/TU71JqaDTJWmIUtEsaT7J6CB
IrZ0+QnuqjALBBCUYQ4W382xn59wl0CAiQPFXxNRh/ARKeNgNt/vDf3X5IZ0TXKD
ebtYtAAD3CMgWQ5xtJRbq3ZeMVuTjsfG2w7r+09zrlZ0jcl8eydZVAXfQ7iLbruF
7f1dPqHy9yqBDhoSObsXlMm9Tw44Ku/NnjuQNP/RMnYG3/NTh5F0qe1969rNBp2U
nCLEO09REnEG4WiGVEZ/QgC431KY4rxPpCi/ZFwEKDC7BLyMWy04DJlutKa16ldE
yxGpph9wDnLFXshrDzmaPK8Xgboz44Idloc3ptYWNZdmb0YzZJxRXUxviFRyxoCp
poi64YoX0F6rHjtHvVJz9CV4/D4uyGOxCkaxYyjQGoVOr10fUfBgS10pHGxEmOp1
OvWb9UqlK8cy/H5ftkNwbqAaGyXt2SztRWBv/YgfMza04C6OhFV2d8K0a5NaRo39
e7+pT0mHqN6sQ7I3r/R3J1FZxWx5pBHn4GZVcVn9/TvfiYooV+ZdAo1e60/RnZml
jaWvevkcXVUhdUPkL5ed/ZIRrKEndXmXQ3472NENvl2CYPQz1iHKCI7py5KpxBvu
kAq3kPlXTrPa++25fgzd4i+qSLU8E3hINzLQDmyg9FN46Wg0OkLYwp66ye8s7Euw
wltbH8e4Fcg96ELUNTPEvi8isrtwr1Ct7EtEMl4fMYU98DzwxQMbgSGD2QKdVTxx
FTQI3OIG4VaOZQetu3jknQ5B7w+O/6pR0PWBAyg8UovtkiDbiqaUCpTAUa49GfXK
q6mquP6i4MrM73knry36Wzyxeoo29Y9IXIX0DRlZUgkeYHl8ziOa/jJNFjpa7UD/
laKtFlsc5jjKShw0Rj/C6cMjbzj66nM6LPnvAxyxDfji4HbPk6JT2QIyWEJT/bdE
xjKdmUGyIzD4j5IjIZOpkTcCTSTB4m8ITQwx8Ce9XJ+t9bkdPfyXPWbQ9bFqv9pG
1Vc0KhVYXzxGMmQVLGL7dcqsYCNN8vjhHg7pOv8z1sIuNTbg+/fsJy8/US53UNBK
CtS2PfPJV1jFJCHfUUze8WW8j3jAK9arSTFpL8FoyykgYrsTda9EMLaSOOG3WNNc
TAPH36TaliUPbxLfhsQJ90RI9yN+jDgUfCyHAxnCmDyVjPmxfP9zaiELa9MJwJSk
C0dHg4EferBqEFQVksbooWnPpqo3g+p6P1ITql8qUa1SMiwMhxlDeIEOqviWT0jg
TNEAjrTgoiusY7RUXQ6Zq+c+2r9A2/9S0kAmcOs8Wj6i+k8Hcv55Vx0PCbZOYMod
dVSogogCKtXkicChF6zDaLqzG2/jHroSQtb4cIyK731EkdyXvdhKlZ8VpZZtr1ca
4ykNjslANkITI+SFBMey0Gy9Y+oxUPKH52d4Sh3ytn1pI8cVRt13f/t+KTHiS274
MeBFcKSnqkiWmxeY/0ijN7awduU4K9SwUP0TdoF4ZzGGK60sz+eVtmKhDIWdi4VJ
xAvTHdIP6FW/2x8FyrywslycxlzWSthyrC3oktanbF0MKIMfaF6bUDgkS/vbe/5N
SOd4eM3L1s8bTXPpRUmXZUNeYEWS98CPhUW/uUijnb1dPIKT0Deh0IRvEKbONB2Q
kYhHRTvxDBb0DiUvdEfJyXUMYE8gfLy5DCt0wNuoE00cb/5E2sOiCTl0WtShzgAy
issowiiAxXAhkT1x4O24iVchgufhm5ieGRBZ8QEuD3XHqQUNgA00GfEDIG9k860R
pZMFcPAamnGgWKRDFKMmuaWO4rdQaf8zC2+3up+35hD3Cr+4zFgB9SUDrV1wvQX/
SbwD1/Jr4DVPcnHFNYK8Vrln+jxakEQ/TJxKdIDklKkqh7FLp8EHqeO+U4QYB3NO
uM+q9qPZYo3Vh+M4yEzrrxPotStlzhjZjg3svOznsvvuKagBtvhRK49WJtnTGqdl
yvw9Ml0BsbYEDJIBFGuvVGrkYRXohQjTZOylz8usWdiVcqMqKgNRiGf2hO4IAdc7
1u1GLoNtLFpdrPbDvxzAOrdtw4xrjUp8fLD7bufJiS5U/voKh6N19uDjc9h0ThLC
G4bxyQ+ZqDQeG6qyKWYneAbQGMVDDgaWJmA2/81R59gF1w6bYGc2dUEjF8jdv00V
bcKUNjnwkmKoMj5JViqOwQYmbslnbdNJqCdBqjlS+irWHCra0AXzqrhlEgG4fFpU
BYyxv2hMM+VpVEN6++6HmQp5hWKxWssLWwBO7b1kcT4qUaNq6+dVI6A5fcDX0Nrz
i0rgMwP2sdWWq2vZPg/NJ9wVHCivQSgYvj2tNtadoH5pysKajtNHG4gnU5tGhqtX
o/akoYj2VcDonaN78ZW8PDRRLCtwvui31U/+bTWZrmJpiaPhMN3z/b2SKnSHQubN
RKXhaiXybfAe0P8i9Qnqo2HdD8/Y4+QHCDQJRIQeuU97auGhZGVTy2rVISAUGdc1
qQa63F2ShQaJ0VlgjTDYreCzZbPHpzewzGpsYAwezyyK+H/ekwTmoWpjpod6hlu/
PiERuwN2kcU9wLt3Gl8NiolqBVHy3So07A/8RJ3Tze2nU699NawCjD7g5nZ3wFFe
TBulpcssQnmDCwGrh1bSWob4Oaes1fPzG4YljLMBbgMh5X4My3dqkSmhORFtkmLV
BlvQNigmviV/7Slz6W184PJo61AORivgFmJbSqLKAVrBfnIs6MwZyA/MJqoHZQRr
XA5CIbAKu99qvQNa/FjlyqjUFLlpNVVg6dtVQoDi6NyzjCVdbt6hDA/3fcvrShu1
+dUAE3zMtqyHPVkGZjwOYaHtXEHkcrbG+Uz0IO/j0HP2Rkhom8/yWQ+5Tsuz+wE3
UjbWQ4Mdo4B1w6aL53LNF2n+iE/ekEvX0n0dKA5dHYGigWbtxjsabetR9F3x/SoB
RvznrxY23/VrZuefBHUuY30a1UnpdMSjC1IYVuGfgg1ZmcQLIGYY+rNeVzeRNma6
ZHbHBaX9AwIW6wlnE6X6XETa9EKx1oMRvPKtJh2O/ZnUudLzlCtDREgBaRfY21wk
SgA9V7D3hYwv07E4Rg8IyPdCKxqSg8linco3ai6gnCVhWh4Y+EF9z6m2BNAN5ipF
XNs0CjVDMii0F4dKoiM1e7wkV45bEKF8Nwc6HhiDTr9C3pNPKWTjJDTCh7U+Opb/
oATBBGc21Waxzm9iIJGGr7p/sl0xMIew4nm3yN+uHfaHMcJ0KB1N/03btBfWIrXy
U67/oHVODBUuCWiwv9sqKHP09wlpISGW56Wswht47YjcRWvbPH6LuZ89oo7E9Rwt
mOBR0jwBal5NIZBLZ0J1hANp9zXVw29FW/Ot5IYXxF+O1K1a4IT6ae18Nds+BxG6
gde5RoPFzpVqKl847iQVLmUFtGyZ6JjF1B6IPr04XPFfLu5zASQXp13aQiMzxZHm
6Mg1gpNhCRxLzwECZ0xrVJvn4brYqXoGFTjXztEYm8VRg7mbBS4Lu8uWy4xDk48S
BK/E5qoVzgEg1FdSlnYVqaik/KummYt8fxVhvOAwXr5oco4hFVVAdsD31nKVSy9h
rbJWAw30EcZBSg/LAH/jUpxRrqyg1rVzBVDNp/9FHtSXHpliLF6cDuM7WRC84wYk
YW+JqRQYH3KroY/6FV8nTgfELuruVR7OI0JGJvqPhlJFT5Kx4VZla2MliIzc2lx5
FABRh4W9F0mZbLTABoTaf14lFIrTl9ALjj0foEOn84hMsbqZG9oc7wwWGKBVxUIr
3DniIGCU8DI2Pv/RVnCaKhLH6HqYvB4NOxszZ2BqwOprd3Y3V/s1sQDVDeTmeMRa
QK0i68vX+s8f+knGtjdq4BJqvNWW98jLmq2kFg4Dk6CnTyu9kvMpbDZ7VvrhWR4i
HoszpVxtxI+m1XvycWWXGiaJgfScq6uRel8XaSdr4qloYQiT2UPxX1uPhiqs/mJk
TBMtPuJM/u5MITxiK536AJQr3Z/+l+xH3K5VPITLeMW37zOhX/fgA66cPDCFLbL9
Zm8o2DYEQ8QYjQrMi2gtsI1N1tMER9259tkp7i8SdTT73KUjKBNH5mf7XyBUC8KG
2PZjF97RoJ/ihrXlH7wGwu0UgZvcNmn7VwnmfWNjtWI6+TELyIGl51KqEySyQxK4
miE2MU1ZxGyycDJmHBlJRJ4JdX1CAuhl6ZZduF1fAotopOT59ZVlMPaj2MpfYjBn
PruQ+KAHUSYoEO9jeSS47uIp698gmiqjAA/6NkdsdXOvYoTuZpORtg5kbqnNgbsq
/66B1218HrrYHezMqbGLmtRtTF0R5jg6T6qiWAfXxXO+gIOUZZndJOivOJl8NyLG
l40v9SszlQ/wzbd1ffnDwjIkZsy8P8VareF9RRtQp73fEvotezMLbQqsxV3Tq21t
cHXTqYFMLBO5kTYCDcjCR5jsaOvWQhJIEFxhd2D9VRsBhgtAhbsASW71FIbrn3s2
hduNU3PqzIuFog48N8vTbR/vGqaHHzk3hzD+EI25zqJfZdDhuRkpQG+W/BlVAdXC
F7LXqfwEh0V07p5/Ek4d68CtZVvZBFyupX7C1a/IRHkBlNikGXcRqWDWSPSMjjvk
xevrDLXezOAX4Ag6erVvY/zj9DzJEo8kh6jOXAHUrYjfMRD+jhX7ep2yD2HYfJV4
Zuom65AEmDEyooD5l9JOWT6OKChBAb4s9VT5h0BiOHFzkHHFueJh0MwVRH6VlWBg
eVd+gLSgHCrK3G6EDtNmiJ+D6DK6knj7pd6OqwYT1tObleemrIdd01ZNpAEAXAT7
rKYEZ4bVNDxpaq9SWwgTlNCqpDKFxA36unSEwZBpa/7FiLeIhzX7ux+0zl7fnFeN
3lsX9QHctKpnxQd10l7jk5mco6dBkmRCAALJ1QzbVGXIfMc1E+J9nth2QF92x/l6
rF+JxtCtyuS9CWfgymt27rqtp9lrA1ih3+ZQUMdYw+wh0YwOy3XJewJSdJMMLxuv
20RR6X0DuIzXVztWfGArU7p2Bs3Zsy1jcwPWiP6v4Br2FM+XzmB4UN6zRTZnCVLu
Jhm5DNVewuPyxI+3XV29JBh48WWPVHZH0x5wQZSCR+ieJJykWebxURXKv96KaGCH
+9FjXC1jDwl5Z/FPqXCt0UbTlmppqdIC1G9PvqnX77NDS/LqZn5htqvUt43tuVC0
rME8X8AdMgbomcJBlkXFc5QuRGQqB6Vn4NFWhvZTVFp+TFwAOFqfKUU7tbukuUMO
s6JuzLaMfPaSxfhXIbHX/FOMwUeMh0SNXah0kiSOaA9n27p6hTpBq9XcSEqWTb3M
ZQ0vXRLs5Ss/6I7o5B+z6MLJxpxf4c31Bp3O2Cxk9N4SruOomRkXxX34wD32P7en
CYbkWXYBIcKPvL6LgyByhhxNac/NPOpRscjprhs4dqDeny5pG1QLQsY8PhdS9wxS
rHwGAt5bCH3IZTqnJQQpfXgkyCJMZ42Y6W+/k4aw9qSGhtNVGhvq7k82VLPfSPRn
f6faEGXgUbwmHdMwU2mG/Mk6X4l7LgbjFpp7I7JcXRXPRWpqQ7L+2C63Szgv8ln2
mcKMkFwD/R3hNr5gmu/fF3OwGXKiJTSe4SojxS2k0AwGpa3Dx5wet8Qjj0Tk/beB
yMhgct/mqVYF4/Wj1n+21K44cNJtMYGxMAfDcbccGrID0TIuc4LFGWdh8BoQnogw
9IcXHBInO/9KYHmUCOPAicR8BqzNBHfIrmO8ZB4lXJEabw9bDAbKAnB+Wy/Rp4Qs
WI5HMx0pH/v4JdwpvWPPC0pKS+xfc3p958xijHeGNWWDL4AnyymoeFUHUj9HGTwq
SJU6amghy8LRDeOGze/PF4YVUBZaG1Ri1wJxR6MIMTlvw0JB3KhqfurK2H7uuF3U
/7dcL2oKW1AAQ5wmZsaWlv+ttbzoKkkXUBNWxcew9SnkccKd7Z688MYUUsNQwQsr
aOfxC1vGjoSwJ4sP2CmwhLjai1TKwN0/nH0Zr8t2EPiZlxZAyd03S/GS4f8VONFZ
9dQboVlx6QG88UWZ4vKMw0UMiOFukT+zRWs4jgFL71NrTCqI8kLQvkHFFLxf6+Kg
1g3FAbmvyf30ajZKMup96uqWo/St8M/MvNkVe2mNpBoXVP5nbhyxOQEjGXqXUKYB
WX0yI4yjN+eHUw00tkjLLFEJgCmX2zUJESIuLLGlbpXszhbtkk33YMN4EHFMrIjH
l2gKd3fGaln4QN3Xc5j/zGvfzfF1qfxuPS0b9i/wO9wudVLLPk5ngW2u42P8gsT/
ntqDHchQZFdcI8hB7CI+IGiy4yhB87YnfNjkHMPLmdljjFmu8ZCXo5D8eswbTmBY
IkS1xABjEFEjM5vk7kTSvfJfU/F4uV4wP1jSXj9FM157vIbaZjO8x1d1yF+SRdXw
w61istNgcbJaT1KSmQquca+LLWl64jlO2mDRhe++GuwvpqF+z5nNyxgEeeBDkPgV
Y4WySwZakTiscussQRqabcbZqzehWuUjUgDh+Epc6oAqzHyxHdC5Fd1vH+ms9Zwb
g34TxxD9pvja4fh3HIicwrr7XLbEzW8BGhCyGHgFOcV50a8HTN8yvmymKh7EYu1r
uYd8GuDHokerfW6x/ygDdTEB0ms2Mtiaccd3Vx2JDNO0Nct6yQuq1fPsHpnXLHzf
mcAuSJGITLgZO4wMbBRkFXvtIZ9iDmuygC4hSSsD8Ly+2IBU0tSvP/sgG8s9pDs+
o2N4eeqpzQvf+TWT9msOyA673pEzvrf0w+8zS4k+VFkaBr4RbQ/ENS6d6bj68xju
hgHoJehGd4wr5VxidIOYNAKZzuc54tsI/EWwbEora2TrDZa9emUHRLEDOKQHz7an
KNVYpHM13WsXU7lrH9YhPxp9/mpw41n40DNQ4yiyl5F1KXJQ3W91B4dfIFcrdHbL
l95EeJEOzNqOJlCmC+AeLhQgHiaAHnIVjMRWcW19M2YMrRPurCLTmnztPe2N3tB3
n5Gf4MUD94UeU7noHzniIybCarD1SCokgObQm0pMAJhT3ap79kOXcqu25gdJoYbF
GqtKjifOkMuVTP/h7H6lW9TwlNV7W/7aCJ6CN/Gr8O/6i01PlmtYX8VgBcn9sdvZ
QHNuENwZx9tZHjzj49WFYVXXz55ZdzWzKOxecRSTDUGP58ZfidLo4gFX4uD0N0Wc
/c+4w8P5V7rr+xEEOkKTMfAMhFemmKtenlIsj+0S6Vyvk2kmTqu3yv/XXFNE2gEl
Q/qLOlI5he4vopJmPvuMDQnK8eUAhq6wyNcKhkG1awkgdreYLRNzUvosKZM/+Xq3
r0bQk2JBhI+59o4JG+L9KMZc15BngL/g4FlWe5wGMryMYScYMIa+jAOc1S7u3L+G
78jhszrn4U9zqJOaLLsiQREjO/deJZ316GnSrGsV3azNXfMyRDGE0VZ/WT/udjUO
XDCwvLLYJuzolYW5ya3jEaK8eHQiPFkP4FTcAwElzbnuHt9sHLsOYOmIT0rFYVbi
oLBm517VKzRj9dxLNG/Gr+6w1qEIHk0Vc54NqYaMdhNfj582AdvlGsqULzGvNjp3
xIl/tM7WeZznjLj/e6Tb+GEMA/M89dhCrgM+IRuYTbGZ+6jtD7vjQlU1/M1xKXGZ
TxWmwYbW9uulLBXjlCUZJ6pBMs1ci9fLLCBRmahuHyKtZP0jXLoGy9nlVWMRVCKH
TYUj5r+2H6kxlJJa16CmIFp1zoOhPDJjl4sBVglI4AzF/y5mCC7//BCeR/xXdV65
dWErF2QewWqyBGyWAYFE69Hf7sLOW4X/JmV31XcpfUmrTZroSmyDcGbuA2xSyC7V
DcrM9XOG+0k5XDl2PmnmPnEcXd3KLTBcsGM0C6/7mWFygnKz2ejfx+XyMISv91PW
4XIIMhb8qUw7qaXevMK6SZzdniDv5EZXqMMhsWlVxh9QIAzf53I+e57eB/VqMGvG
+z5z2Z7Z60vO71uW+bgi8uiEuKTwWWpA+BzAT7l4FraCMpNFklFAR9JjcoECIW4Y
PktyGnGLXUMK1Xu411DZpF9uZSutw3NZdLIZxK9LGtDIUNIAYs31HDHmGlpxF5vx
ZLJc1pBRiC687ERx+d3VouR91hyokEL3NEgp+BQys1010RP9Lusqi/r5OvJjYVIX
NZ1URh1AXRSQjjPqwa1aFwRIyf+TMhX0IOsb+AP9BfiVPdw+jslLWftMcnwmtWsu
cnR+xK9mR+anJNDceHAHrDPak6gAJW6iIRqt+FB5qA2fu9abvCo1KZdhW6l0g8Vo
nJPfTQe80KZIda7eHKkH3s1mijPids6KUAJcMv7Ld5RxIvUSzYD8WNwDuCG+AdBR
d1pOx/mlRYb9FTkdt0Io7AA4o6X3ueHbVp2M2063mGP48GfPtB6SpvqEzfXBHGS3
0+Pi4Hp6CvvFQp+HBC+MFcTM/l4NnpsrXYPdViYPo7WTxtQJHoSL0dHVes1tgNTF
SwNpSeXw3lL/aPWohWwopbHxYrUKuaqHG5WifyEI3GQru1JTTeU3ryfO34pWfMlx
R3qrizZ+himFkuavjnbPtMfnfOqXAUKHv3AY46g12b9o3+nwTX4d6aydUIzRg+Ro
pDZLUhIzeqlK9K9Oxm2rhcSLcKA5UI023ALzoikzOUSO+UR0iRncrhnfcp2y8zQu
mhTVtvmCQATT6bZxF/hAvr/9t32b9ImudsWZn9MXcLU2qlrK8yLUPXmxkYm9qbTi
n5GJpcneSS1n14cz/SMGqZkQt9EfqRbiDvB9M4rMDGLx0+BSisZO9Xh7YJdfrriy
pjuUo9F7p6AkQ8DvTZBaGvpuXqwMyMpmjDWwLa/aqXd4SzWen6tP1pszPGzhpxqV
LeZu9eRTb7umV37oeaDzClqasSElrtgcQ1TdEqkLIqq1cE9S8oplsTfsOEl95z6n
18M7d89Uuvmtal9emIcSywb4c8wTn0Ie7fxsEDb/SjZwjNwwdXf/cOX6AK4CrQzl
ybWAFi+mmGxmR6j3itUn09AFadGXDSnLHNdUPL2C5msRf8uz8lC21u5+NBOmRjwF
/TCtehs7nbb0+ZcmeM1SKbbEdWA9tZc0UQOAkgF0YEYXDkE+WgZZwnu8DuLuJ6PV
p5d9ZmquhBgT74Ws89mWKfhLUpLci7CrOINXMBVBac1Zqp5YEy0MSYvGF9akz4XL
zraShf9SnGbsWdINd3JBq/98+Ieq04p9p/F1rarDy3wBJ9VcYnD6cKE70yS3vdj/
lx3hoFKj1vEGGo69PjKKBqu9+K6IskQc/uqfsLC8IvPhUJh6aPfvp1esrq2oeUDN
0NLWBhBecQsaR+7ZQUXoQEqxExBRXJfBrCwX9O6ZoTQCIrH2rme+PPLUuOfxRnaf
6DeqVr3Y6MJNHaSawD6SWt8O2/WDNLxUwDVnbKTVclkr0lpvMDoqA4Nl0jzMYO0U
m03B+bdZmhfcu0+ph+AMkrvV76SYnZwkAeehXx+SGdHY99XiTZTWyEWMZLdoku3b
XgSQEi0EymOCtr7fgEMDlZH6BwWnTLmXcK5RUVgcs5Q5dYUlXCcGrUZs7B78u0Nw
ie3APf9OlurCHMSfT7TwT4vKicEgIbpS8mEbxQVA/j8wgf8/Objm8jr2EE1F9VhN
upowyr5dXUzteuHsApCjMT063ASxOAD9i/0rpNJzmlLY5PrkcSc/OxNUZVSdMRB+
Db8/nPhxuSZJbG9R4Q+DcdqHzAUQwZglRUaLB7wABqiv4XT9ojPzCQQuBBhN2Qfw
p3lX/I8sG9VgfuEAo07PINC7jy6sWFrYTKyEgnhtspKcJC/ljbiiskn2rQLsvSIs
db3cuNH5Eb2+flk5mgPqJjRPmeV3o6VcixNLzVO30VlNuFuIcR1nxVTrp9g4hkmH
r6JvuSvyw2nHrldrNPjHUaqTdzVXG6oHwmC4TDyFxs782iZEqqaH1trfz5yOdIjK
drw827jNAmSDPNIW8i2wPkqCcBwortljkMrtW+ZPSLTByaQ5VHxyVgq+dGfdeKR7
M4e+mmmmDE4tFIepYhFyVX5ummDkoMzeHuZajBAg2Lz9EpUITPAxibjyko9Zfr+5
+5xjnlN4MClkq2C3s5Qg+3XMw+GSuqjd7OCkkbl6+R3HSLUABOsEDKI6ti87sSEe
PgEoXC6a2lVbinCcCUk7XxiuxBtEy/ISwG3uy5F6ZhlY7HdidOsLNcJYNXCa/Udo
PY1sM2zJAnpBzVfCtpDi51BVoDYowTrZkp4mElwuKxxfonWBBplDEryt/VVbnboC
NHBXUNQQh1tCqp/ognBvE/gQz0AYUH8shqb6klOI4kB4Rlrt3Cij29ncK1FwnqDl
nQvGEHp60FLSfHCC0f354az5W71s7o4wfjUVyJpV5NKIGuhfeGBTLKURLa5GJAJX
iuhHGZ7/+jJrBf3DZRCZmHWuswnabHcFoCLh6udvDx3ZHwMU7ngEBDMPTepZNyRJ
1DTOVG1U3HjtGFSgE0G8NcVo8Da2pS8/nEOeQVnf+rloW8ZxX6Kv9jR1rCQGvQEc
jIJXHMiWKnEy96qXcWKzs94f9AgzdYoGsAoRfMMFNFaLyqM4VCHjCrKqYFBvX4gH
C/4sNd3GaHxsoWkZ5AHaCADT3T6TC05lhLRlug4O4pc5HhoiWQQn6K3RPGjShREV
kQGkrZ2MCJ/SupQcuMyWP7B2U5oY3VT5evOMO784L3s4RpfyTfZ2qEPgVb88M2Vj
w/lkFIqTuVuyGBlPCK3p1FnHE4FZhtnCYFF2o1MAKCk178de+8ArXMXAgXJy9k+i
P2uVRBkf/qqDjPfDrH4Ju42P54XpErxX04z9u0+NSjJGPayS9MO5NuHEzSMN//mK
aXXX81Jhto7FnQCcon1TF4WsT6f+AWxMGHSXyTj485cov0UY1sSWBk1Amf0nhAmt
VXI5EinTu+D8A5jEF7ed97A/GUcuS5k16Trixntxy8evMyGSpED5Jt4vm/Fv7J3I
44CtaeqC+VUPUWqfEXsVuiVRH8Rla1NI/nztyCoq0cFJZYH60B2GR0j5fBzAJBxA
0t+o5PycgIYXz1F4Js5EXH1k235/fbZ9BuOKJRIEDEg8JL4APEsrYcVkJELwM7PH
u0DlCFpJA3wvdMohBkwLBsEGlnyAg0wX/7G/wTQihNJXDDdHbHjlITkgtZhHo7NE
Uq0aPyOiJ2Ea4BGq7BPY3lOnp+ahes/sRJXvddY24K8x3k2jvpckO0/X8F/Atm0U
n1KIVrKwodOxgX70QY5v6TqgnJbT3DZYeuMVDTRzjW4WvVmqlmLokzkofqg2Bs3c
ur1EBr7XUPfpRkr3AmdxGLAdGsohPVJMGEnRe2A4HvH2/Vkxanu/YmhlvAveWWwH
M77+U/AsztqQJ4tPB5u93CbWfJzUvPfn0wStcUJ7HAFpaThkKTOJq9w+FIrwaymo
45KK3tUtOVYIZhrJzG2RoR85GkOwPg54tuvDrGkw/m034OfRdqncgEA+MwGaLJdj
lWkhO/YmN5KzlQzistwqgrDGmi3E4ZxYuRw4T2sDXrA9x3cPEghhjI5QU0kk7wXJ
jnfmpxt2yHDiQl9ePacghTR+TI9lbLfkwkyyMUqtcD9Ci4QqU9cem+G8an2ZlfLT
hWDiVZjRN8KYsL6Ym/iFxCUANOC2wUxjG3cSgl3lQQ6mWaUwc46Own9jqW//bOo3
ztwd35qiok3qvLkNeLeqHuo9SjNMMLy+MR4G3TxuAyO4vGP9I1nATWsNqW5JfPpa
Uugkd/EOEAc9zx4HQcuDW/7fjDxSrR1UTzgchfhs+AQVhxZOopBo59nzbBAac4IN
v+NoX/JamNhgCbWAsOwXsQX8ZhPJzFkfL7MqL20uDHdo7Sme6RoS/x0pgtrl0Om/
325bnQAoZeHSD+l9aJcdbTdHigh+/Mdasrs1ExA9I3YP/BotaZjhp5K+uWlHqXRU
R6ocMIFAsjRuTphPQbpGXLeAfk1xBsHHl+pRerSLzwR9EcKrTNidXClgLGEt8YLz
xmSWECYwm/qfW3voOBH3OSHjxSS/L3No2U5IdYYNMl8JnO2Pe8FwxftZuuOvf/C2
wRYsOH0I3rouvE4ju61Rb1mtxSNy7KeS4L2i6nhf6iBmqYM8OqAZKni2UHxgKjTa
Rml9IwddsmNV1CPR15kiAnPyLvS85pXFeAfOvDTrTQxuEM4kBZwK8yclGg1fumYr
SykGdxGCrq/r+hiwD+nYacfUkD4WwWP/xJkQlHzqtP+w+0SqvgOvSv2LPV4rheJZ
gl5fYgi+tkMB692a8DxzHTSpsVXhr3czXxhhfxA7fFK1UxkfUKdquknPkRbAsfdV
E4JOpZlnCAHRC9j3cvnOzWQS0NKfH2qafX3zNv/rv853Brv9TIUcY8voH5hXhDjC
DQaYAUpt9KskXAQwK33KgyQX2gEXrFvSjSBsNSeLJ1GLmFKHebd0WFc0VcO2Nzt0
yPRpDeU9Do3zKdh15ODLtzI3nXTTokhg5vlQ7Ci+ZTU=
`pragma protect end_protected
