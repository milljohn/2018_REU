// hps_emac.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module hps_emac (
		input  wire        read,               //   avalon_slave.read
		input  wire        write,              //               .write
		input  wire [31:0] writedata,          //               .writedata
		output wire [31:0] readdata,           //               .readdata
		input  wire        addr,               //               .address
		input  wire [7:0]  phy_txd_o,          //           emac.phy_txd_o
		input  wire        phy_txen_o,         //               .phy_txen_o
		input  wire        phy_txer_o,         //               .phy_txer_o
		input  wire        mdo_o,              //               .gmii_mdo_o
		input  wire        mdo_o_e,            //               .gmii_mdo_o_e
		input  wire        ptp_pps_o,          //               .ptp_pps_o
		output wire        phy_rxdv_i,         //               .phy_rxdv_i
		output wire        phy_rxer_i,         //               .phy_rxer_i
		output wire [7:0]  phy_rxd_i,          //               .phy_rxd_i
		output wire        phy_col_i,          //               .phy_col_i
		output wire        phy_crs_i,          //               .phy_crs_i
		output wire        mdi_i,              //               .gmii_mdi_i
		output wire        ptp_aux_ts_trig_i,  //               .ptp_aux_ts_trig_i
		input  wire        phy_txclk_o,        //   emac_gtx_clk.clk
		output wire        clk_rx_i,           // emac_rx_clk_in.clk
		input  wire        rst_rx_n_o,         //  emac_rx_reset.reset_n
		output wire        clk_tx_i,           // emac_tx_clk_in.clk
		input  wire        rst_tx_n_o,         //  emac_tx_reset.reset_n
		input  wire        mac_tx_clk_i,       //       hps_gmii.phy_tx_clk_i
		input  wire        mac_rx_clk,         //               .phy_rx_clk_i
		input  wire        mac_rxdv,           //               .phy_rxdv_i
		input  wire        mac_rxer,           //               .phy_rxer_i
		input  wire [7:0]  mac_rxd,            //               .phy_rxd_i
		input  wire        mac_col,            //               .phy_col_i
		input  wire        mac_crs,            //               .phy_crs_i
		output wire        mac_tx_clk_o,       //               .phy_tx_clk_o
		output wire        mac_rst_tx_n,       //               .rst_tx_n
		output wire        mac_rst_rx_n,       //               .rst_rx_n
		output wire [7:0]  mac_txd,            //               .phy_txd_o
		output wire        mac_txen,           //               .phy_txen_o
		output wire        mac_txer,           //               .phy_txer_o
		output wire [1:0]  mac_speed,          //               .phy_mac_speed_o
		input  wire        mdi_in,             //           mdio.gmii_mdi_i
		output wire        mdo_out,            //               .gmii_mdo_o
		output wire        mdo_out_en,         //               .gmii_mdo_o_e
		input  wire        clk,                //     peri_clock.clk
		input  wire        rst_n,              //     peri_reset.reset_n
		input  wire        ptp_aux_ts_trig_in, //            ptp.ptp_aux_ts_trig_i
		output wire        ptp_pps_out         //               .ptp_pps_o
	);

	altera_hps_emac_interface_splitter #(
		.MAC_SPEED_CSR_ENABLE (1)
	) hps_emac_interface_splitter_0 (
		.phy_txclk_o        (phy_txclk_o),        //   emac_gtx_clk.clk
		.clk_tx_i           (clk_tx_i),           // emac_tx_clk_in.clk
		.clk_rx_i           (clk_rx_i),           // emac_rx_clk_in.clk
		.rst_tx_n_o         (rst_tx_n_o),         //  emac_tx_reset.reset_n
		.rst_rx_n_o         (rst_rx_n_o),         //  emac_rx_reset.reset_n
		.mac_tx_clk_i       (mac_tx_clk_i),       //       hps_gmii.phy_tx_clk_i
		.mac_rx_clk         (mac_rx_clk),         //               .phy_rx_clk_i
		.mac_rxdv           (mac_rxdv),           //               .phy_rxdv_i
		.mac_rxer           (mac_rxer),           //               .phy_rxer_i
		.mac_rxd            (mac_rxd),            //               .phy_rxd_i
		.mac_col            (mac_col),            //               .phy_col_i
		.mac_crs            (mac_crs),            //               .phy_crs_i
		.mac_tx_clk_o       (mac_tx_clk_o),       //               .phy_tx_clk_o
		.mac_rst_tx_n       (mac_rst_tx_n),       //               .rst_tx_n
		.mac_rst_rx_n       (mac_rst_rx_n),       //               .rst_rx_n
		.mac_txd            (mac_txd),            //               .phy_txd_o
		.mac_txen           (mac_txen),           //               .phy_txen_o
		.mac_txer           (mac_txer),           //               .phy_txer_o
		.mac_speed          (mac_speed),          //               .phy_mac_speed_o
		.mdi_in             (mdi_in),             //           mdio.gmii_mdi_i
		.mdo_out            (mdo_out),            //               .gmii_mdo_o
		.mdo_out_en         (mdo_out_en),         //               .gmii_mdo_o_e
		.clk                (clk),                //     peri_clock.clk
		.rst_n              (rst_n),              //     peri_reset.reset_n
		.read               (read),               //   avalon_slave.read
		.write              (write),              //               .write
		.writedata          (writedata),          //               .writedata
		.readdata           (readdata),           //               .readdata
		.addr               (addr),               //               .address
		.phy_txd_o          (phy_txd_o),          //           emac.phy_txd_o
		.phy_txen_o         (phy_txen_o),         //               .phy_txen_o
		.phy_txer_o         (phy_txer_o),         //               .phy_txer_o
		.mdo_o              (mdo_o),              //               .gmii_mdo_o
		.mdo_o_e            (mdo_o_e),            //               .gmii_mdo_o_e
		.ptp_pps_o          (ptp_pps_o),          //               .ptp_pps_o
		.phy_rxdv_i         (phy_rxdv_i),         //               .phy_rxdv_i
		.phy_rxer_i         (phy_rxer_i),         //               .phy_rxer_i
		.phy_rxd_i          (phy_rxd_i),          //               .phy_rxd_i
		.phy_col_i          (phy_col_i),          //               .phy_col_i
		.phy_crs_i          (phy_crs_i),          //               .phy_crs_i
		.mdi_i              (mdi_i),              //               .gmii_mdi_i
		.ptp_aux_ts_trig_i  (ptp_aux_ts_trig_i),  //               .ptp_aux_ts_trig_i
		.ptp_aux_ts_trig_in (ptp_aux_ts_trig_in), //            ptp.ptp_aux_ts_trig_i
		.ptp_pps_out        (ptp_pps_out),        //               .ptp_pps_o
		.phy_mac_speed_o    (2'b00),              //    (terminated)
		.ptp_tstmp_data     (1'b0),               //    (terminated)
		.ptp_tstmp_en       (1'b0)                //    (terminated)
	);

endmodule
