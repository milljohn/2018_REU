// adc.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module adc (
		input  wire        slave_clk,          //     clock_sink.clk
		input  wire        adc_clk,            // clock_sink_adc.clk
		output wire        ADC_CONVST,         //    conduit_end.CONVST
		output wire        ADC_SCK,            //               .SCK
		output wire        ADC_SDI,            //               .SDI
		input  wire        ADC_SDO,            //               .SDO
		input  wire        slave_reset_n,      //     reset_sink.reset_n
		input  wire        slave_chipselect_n, //          slave.chipselect_n
		input  wire        slave_read_n,       //               .read_n
		output wire [15:0] slave_readdata,     //               .readdata
		input  wire        slave_addr,         //               .address
		input  wire        slave_wrtie_n,      //               .write_n
		input  wire [15:0] slave_wriredata     //               .writedata
	);

	adc_ltc2308_fifo adc_ltc2308_0 (
		.slave_chipselect_n (slave_chipselect_n), //          slave.chipselect_n
		.slave_read_n       (slave_read_n),       //               .read_n
		.slave_readdata     (slave_readdata),     //               .readdata
		.slave_addr         (slave_addr),         //               .address
		.slave_wrtie_n      (slave_wrtie_n),      //               .write_n
		.slave_wriredata    (slave_wriredata),    //               .writedata
		.ADC_CONVST         (ADC_CONVST),         //    conduit_end.export
		.ADC_SCK            (ADC_SCK),            //               .export
		.ADC_SDI            (ADC_SDI),            //               .export
		.ADC_SDO            (ADC_SDO),            //               .export
		.slave_reset_n      (slave_reset_n),      //     reset_sink.reset_n
		.slave_clk          (slave_clk),          //     clock_sink.clk
		.adc_clk            (adc_clk)             // clock_sink_adc.clk
	);

endmodule
