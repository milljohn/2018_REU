// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0.1
// ALTERA_TIMESTAMP:Thu Jun  4 11:11:15 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PBxLvGBsXMAD/FcwbAOceb0CmRA9Py8GUYkdl+NqUcl+gBmpDiv9+23NVmb6rS3c
bob+m07Q7ouVAFvHR+nnbstvZKLwMTtNO3EsSD8w8ArVlhiJVe7PF8H1PLFza1Vo
iiKZBvNRTHisJjc1rHgWyQ66w+xR2AHYxljJsKshR34=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37216)
83DYMeBlRtOH7yd4dCLR5Jkd4kOZHZ0d+EnFHQs3fykvSS2OmOhI4HGHJfixKJpE
kpYFYJlWHvckZfhluT6n342LZRIhdbJxDRz+MsDoNJ92xjOHa/WGbPAL83ZVOalr
rrwvO1YfSDcuAhZuw+Z4zwPnZRAVG+g27ekdg5pXfzxh8rX4I4aL7RxLPV/6lmS8
YGBFL5lm/teb+dr1q8ecR1QFK5XJc30d2Y0TlNrpO6alcp+wAQZMClh3wYkmCpc6
RSBuqJ3QRyyLdtZvtlcPcJVkl9/ERe4uw0X5WNDqU8QG4NKgQwEYhSqWNW6ieDT5
V2j9+j4ys8kcuvZXGk+x+pghAQc5zvuQRgfwwrLUyzY0W/W2tINDAnTNIu+/nsAm
sve3p6PPU7zIZIwh4rvGAkKeCSuZv/ZP3zi/9bWcGpVTseGb+UJ5on44LY54VJxm
y+xamBKhsmgQzJBr7ZPlJlKZlo2owHTbTFk0LVvsLI3SW7P23cGoRJ1sHzuUiCKU
0IVocmdfpCQpuO6sXVjIj8I/IcnsK3dmjnLKG3yEbe4fAsQQOqHZoi/9M6izfQGL
f+bPtSFA5X6tl1VWuy9iee1VtjRtbfAkD6F8laMLti5H2MwhQ9VzjOY2NRTXarH9
HGFWsIq31YzML2VqYlGjkg0xM9iDHCC5GYgze5tcEfh4cRs5KQV1hYgqRfrvpi+g
valesRDbAVkJkxxebtvGNkXaurhailgBDRHSKuPnpYcMkQnMTGxzqk6+bO8KzAhs
WNl3XKGJu7DSxYYHYsMXIm2BB1FAxb9bxLD4HpclVx+jTBYHhr1ZxYq6gYgVlE2y
G102lqfXWj5f9elAqzeaeo9fWAdUWu//tQtnutHfWKKwBKOkDA3Ge7sQvvFtuIHl
vlfaVJKyn8zTTKRj/DhetESJlMhHCnHnX8QoXiuGwRzeld6ZX+39CuVFQTviUrqu
TWIdEsEo/v0tM9rTDvJNCAzna0ww8VXEzmBRZmx8Is+uapSSk5uaRJZfptMLqPZ1
8nsYGdFBnoU2Pa8jfnBSyyz8msNwK9U5AcRkM6Fi2fZFfzCttx91LzT72pcGjqQw
bTzRl0yCe43sgJyjGSW7b/FY+5d5WPP9F1V4pImgJeKRF20lyf/KRK9FpLMJqIX5
3R6ph4oaWAZrz8zfR1At6ZbXSPiN8nzaN02r3WVaud/TlCB2MEshDgxGP5isKoWN
K5wf1kna8Udbpyh1Y99uHm9brVcfDpMcL0/sfb2xm5BqGwiXnV0RN+0kSef6V4fE
iE1KnHRXyzXwOOKqN9iiOjqNGq2nRCf9PlqG1rF3jckO0QSThfdSx7cA93KUYND/
YNmQtXHdRUUOaMwp8i67cARioFdceHcQFcczw9VUhSM3FOAPxHMv0oMuY1vj3kGj
K2rDnQkSGvmjaBpdfwOBSWfFYBEDRyZW4EjhEp6Ux1q3k9txXEQyopikLcyNPqXR
njcEsrKKtrCp26caMCUTv0cU0MTfDACRUErGiFkzD1Jx2hHeTBfSDOdnPFrqOqzd
3k7FLn6UcTR3MPS1nLxiIBkv61NUkbAUa6Dr1y1lGhXEx5S5h6ZFChO+WKmpO4Na
uhRrLBT/R+fPSfYq0Vt44/GpVIqMyEPQrwy8JHO+PpPe/MHE57NnkDtXRN36dGaK
5a1fTwdWtoVjgQFZ8clQZ2MReBpMto36jhF5+nbRix1ErNvrXwEY72ENW7lBG7LR
DlMRz6hxd31F8VU1N9ILO7ZHTJUqIQlm4GJNbjF3dkBPV10tQZWVy5h81YN27AzO
WMbaecFzaRA8sMFbcC7j6c6OulTEwgpOX00IixFfDc4w4cENNiyyntsf7ggAKO5H
Way/YTA2OfuXB7AflPaKMK41M4DBhrVW983dyruwbZRA2b83+sMiXdR4u2LCuqxl
H75ytlmAW3th1QhNSWEZo9CQL4TcHbgT/YjFzGiTzEZXdduqHgg11zlSpiqwb0Rj
yLAXhNC6sr8XINQQQEotGaXy6J/bxXWBHOePpZ2Imas8KDkYZ+TwY+bxZiyGnZOi
4W29N0VKWdbsOKFYwdgAxU9gINxBpBIasapa87Qn7CmTnQ7fjBNlmNlq6CkZ3Uj4
wckYi9MptivIE6Be1FhPZBBj1A4Dx8JR/jgHHk03p54b/Tv9k/JxnjuWk0HFfSf2
G8L6NQJk2Y9OF1aZE2Jdk92vl/oO2ukYUi0z2vv//4zHwL3QwDgReWXYfJ0GCnUM
4mNiVRu7NzA/rJFHDRqFtLeQKXVDGO89oHKVg7ywL0EGSRfbwz26t4fQIFBrPJPF
DQc+001PP+Zk7zeTYBWW8p/HlKjyxBOvVBnWAWvIMFnfHGUYeArPdNXMxXZqZ776
Wi+Ak5xZgIXy6JXUQ3KU21Z55UmZhg/MFcSya5mrNplOBzWwT9EREttHNjwiZZ0M
2ctR9VwJygqCL6Rnfilb+m8iEK/SLMgK0ItcVGjiCfpDy3SanTEGIdFGtI0vQAOI
Za36GriFOi14siQ2VZQZcgR9kZL+VjtFl+usF2+sUkLsv0iNJOSmn8LFH7mxWkO7
L44im9s6H0BIgFN1Q+LAjoUlh/6eYDvV/LQBeSB6SDPtHGayhuoLpPOgVkzyF7qo
2yfxv81aEyoUwKfI5UQZyYHx6QvTbzMMKMB0UohWWkHk2LoIQV8ccelYOOl1pmTN
vX++YpPrgNThJiUMh9+g1MoSYJNxomAJkDC44HN6sd2Rwq3V+bMeJiBBwwqM+hQD
jCPFLHTvMR7SamuzUwVGWTk2IuqeyO1YOh7JGreOYbbyfl8dtpX6FswMglSaKgAB
5Zq2wLukSeoeBui6pCKXXSDEYPPw6pX54t4Ogh5W0XyobOlAEgRYtd4rCrZjitc7
koaFl7AeP2JJ5oZNI3aicfhhRMEXTV9E29j9ZrHhdf3z2oRcKgoWcVcZ4jmWP5Ws
n22zgrAHBOF+fMJrcUHy1w4lQ7MwI085Ai73yAAmVpeCPLA10ZHbh8QH1iWPbeoA
6IAVZ3lf19KK05uqSjETEhj+/excbkDvExfBFyHw1GPa/N+s5wASTWLaiYT+51IS
Ore6HFcd5BbLH4G1jKOooJi013p34uG4apqciwszS6why7I1rRZWD5+I7XAFS6FQ
Ebf1vSwykugM0LL/RiRH06cnC0HtzrPSw/ccujQP3Bl1pa/gbHLPPaXPi/g61eW7
jRwIMmm5UFUOS/bZh6ikGaCjdJdtZhCA/UHwD1gSGpF5Q6sbDSqpgLu1ADx0RM9X
5t5yEPMxQuOB20bw64fNKFbxBUuhxOIdnc5ZcWzjYh0DooJaJuW7Yg8OIlfj7Gfe
ABTYKE7krqzW5m/i4iw7suad16/j5/1MY7HDBKxs/UHEEh+ohu/YhKlikN854t6k
sz9sinzYBnpCt0U2T5Y+QPP6/qwIXRy+Lp2X6xTf4n0HJajxtBoYrWu7xy+0pQgR
/u/rZPGC6WICAKAGIGrS6scCMl42WRWrGlqpddQQ/EdQakepka59W0toVTEmOBXE
HZm4tUUFAe5d0taVNTwDnNq2bK2AJWw6MhzzZHdIfP54gDr6w/qPSMJc6iVxRinl
xUBLlhc/XcxuWYPooRYc5bpJWOVYLOB498RbRMXfTB631RtL5tIXaoKipEBJ/Tk0
pK38yrNk2ODJxVEWZvj29wzirXHPNF7/gNT+YIeb+WOYo7HkTpTH7ih7LK56Md5d
U8y7zRPdNpUELmPAc35LxD/Zf1Q4r1SKoMf+vdiOASeyR2k2G5ua6FKfM1pUDH0J
2N8b9fP/Uvxc1qUmIwO/VLB+8eMQ/Ys/Wz34NFOZdnO9hlIGEHMF206FRgw2sA2M
Xk+XNiBS7U0d93uSX97Bj/pZWD7pQd8+M+Ti9fV0F4Kl+JkyCQQhfJp52tfxhrPQ
/t6BZKn62qf9zk/0S+6eoSVaE06TFtguzQnW9a5y6CbBm+8vH2qKQ08moioCHa4y
KzqGXxQJSJMtkXWnk8A1UZ1IhmiIUGSoA2sYPmXb9Q+JFk3dGGj3wCI844f+RMZO
GLxFpCwxxQ/+85n/uszEn/iSC1Z77kggKmtFcraPQRJkYdNilMyodVcdC0ancqrP
D8fPnmVKEba+4Px5gEyaHL+PwvFYTQ6fuu5dbU+Hf9oI4418ego04KYXo3ISfRuN
QmtT/ZexTbPdyqgDd9siL2QsfZvKvQzYls/8cpJKUlwZvGWuMtyYfmyWumQCOaPI
R2M6tdkKAFVeg8o20uii5mlAhdzTQWCsIyWHLoEZDty/ZAO8SvZVpnfPiyCwa/WC
4I426xG25Niwqt6q6HP4MMGjgQVZeLYihlWjl6pI1mUPY4+ZwqHh4moifawoXjB/
8fhV+4dsr2YAPSeZ4V3TzJwXWbaIrgsKApXBsUWq/+zfoP8iXLkBBZ5WHDp9oBZV
6VxAY6AACHPHTwVIJVDflCukXurXnhkCYvvnyGl3Hp08vAFmgXk6UTnTyzduhBFC
4ugcUOQzOOL68+oDf8iPwOEFxIqLhTuc0IudjKMTEynQKiU9vJ74qYrAak0HFT/2
LFKD/+MTZajR3aff94tbaHdBwMWig6+edHre4TmCWJiKMmtJpUuhQfbz1Ejwrzjc
NoKaLP3TbucW6/5/wXOTxpg+VJ6BFktuYy4gPdS3l5UY4rSrXm/uzL0kMx63nNIJ
eDfCIaWD8B28NvSKxkIbAUDalhNtdPKiQBKKzJoamEk7017zIJUQe5HLDH2uAzAf
dvcu1TcnLe5ddFVDTBvGcihz/52SWd4kPHws6RTXQiH/aK8kn2lNz37RCT502ioM
X4bPURHCcO3M8U/W3sqcqlv3vpNawRXZuOw6nQb0twfyS5n3TmOsOz1L7MY+tYo2
n60KdGBeFOae5c4A9IrzgAf68Ph7EGewOTBGFmS0LdZIG7QfsVwnD62KOzIIUj1g
0CLUdMZphaTDCv1zGZQLoKUtdSdmUVgui1G3VxnayPNW+xRtWqPc/ijJRhDfxlAr
G320KZWSg5LpTe53p/p0sOdUdSmBWKFFABuQpBDh87aib5V6EHw0WDDwleDIKa7x
S8dzmlHraqrT+faTlgbxsu6kbygZBCqPquRC+jQA71TExRt1QJTIw0SfWOCNT8fG
RvWQG7tVulYXDG5V/G9ujg/PsVd3q1uJxLlrvBRbrowNIxoxJ5mLsZ/i7nRJqWPw
l7VE0slo4M6bcAfVB0z5WL6QWlnQrXcIfKaTY4niX/OXhSDQqGH4BZO1dBoaYWFC
cWWUBNWKSxdMx1JAFBFo422iGXXiLz1qyslIKBcDUBo1DZb7cd9QkRkSCuLXW5Zl
CZfN3tW6cDa2uLVriqL0Fea4jgP4W3QmBlMNwXtmeomHVkGWNTwClQDjbYjGt6e+
D0ZvggdQLq6z37u70IU7TjbYjmK+itO2uMD2G/Hsb8LeEnLA6UOSbA3NkJ9gNjGo
1mBv+FjmOR1/q7G+mw34Qcy8a+A3S3xs/qecgyksDa87j+IM2bSwXybjCY7RTyd9
Ayksimgtjp/UIS422yH0o43a6tuRF73JK7LEeQBzZ0iuwB4akxyLc5F1mZaxG1VA
zcwWyL8UGfhATaSSSHRXlhL4OC+Y/w8iCmljq1M1RhOVu66rZ13doa0etiirq90w
rN/sSNbtF70TA1fGyoIdQkcvz1JAOw2cXeMZBc/j5pf5f2Ln38um5JakDkM0VBDm
9BKJk5h0Ws3jWe18HzYQys0QeNzBtqa+gv1NxImhgRenrFIUKvzHivYEQJN5fB5G
rhjfzetWKjOh3rYoeK6eK7/1Hkw+j4RKz60OfwZT7edz8OY+QSdYabKnXp8fa5cR
yEHIodLqRnD/clxuOcUP8W77Fs0EXhkgPkQFMWqXAW3v1KdHe9ftTPOC6zZdPWte
TEBQch3W6HINmTMGYalwSJ8NuI9IHinVpOq9Wvb+DGHOtQpeLK2dyNkdHw3x/eEk
Kn1KjIOx4gJwp3UifY1gPjOazguAr5dIQGl0UDQOEcabIDevSfVjgSv5hzTIl9Kh
oICBYjFkdhDjKOVY1fOxZdhgzLe4JiumMoa+p9i8G1on/y0RQvjZ7lGQunS/WkfY
5Cm8LFMcvwebuij+ZbDoT8UuCO5I0XE5xeajqz5QZr8E/LXTIWuAwxL80isJBra1
vlfVdEQ7pztuhE86Nb0jkwz3gucDYyx54Q8BeTN8uePLXZJBnnj+m5wQ/ahpV4P5
sMGNGCiMKAnTj+5aIjmiNj04twyGwLpU5Htr8o4ZpKemGF/y0uNEj6S4gCGuKY8D
xC9LC2xQzrKK39qgOZZIhX+UJFt7kAcKfKcfhkS/bYhniU9uCQbb9jECEqUvIQMi
eYc5HT06d24BT/Sg3/IWv54rTbVALF5fEum3w6JLb1eZSUcvRlQqHwGpiJJ6XLH2
lD4Cy+DiGw6UomewqedOoPwQQ98uY8tbt+w5iwp19vyvd5ex9roEXj92e+1CRfyF
6k1NyAu+DoICIf0E1SotEYcpdCAMCQDSy0dlxwlLVBfR2iCyA8zOtqAThAH9aSYJ
+DxF/3432ocWtB0ibohFYlPVed0YnCupIXqu+DpACoZGP+gq2RnlK56SdzUSHzGU
IhqOfoJ1L7666GwAQCE8anqTBF8lY+xKnQV4+L21AfDBuBvdkc+PO00K8ol+TWK+
dJDgb5FkDSRAMZWfca1tTDzkRZ2bMSQYor7FqqzlMscpjMHG8ZH+5+ml8v/4tD6J
AmZEz7dVPEyzYI+so3jyROtUa3NBekDVtoJwEUfYpRkUMxxc9FxWCkS51dowcd5a
g16VazbW8uq3rxpSWp2jQEx9FCIxlT/xAIQ2lSKL2jvv2Uy07UWJRMRsKkmAkwDS
qQeL5v+KuQ/GPjobb49tQ9NUsh2kqsK9cX/xeEBViLCZ4mSS1v7P8oSGv6vBP7fL
jDrOmABhaWoLCEE2Lv+JF5hu+GrWbBv2vsLxl1SLoztXikJRzgg2RL033wdE1++M
Fj1tdQW0CxYgbMPxDSKmBhYqgQH6zvfbJ4PsDj39xvQ5w+hTWJzhB7iFGynWr90n
TRz2l8GcSvUHvWPIaCjSebGJ5OFCp9F9TQXnBBr9ZTZY3CqFDL+Ti5JsxF2frirL
19aHWBttpXbu0yp31X44v+FedIcNkNPj8l4j3VjMQXJH98ZVS1fkcBwqqBI57rXY
pnzBBbqkRc18CvibV91rtk7lEJnwuHVfjdtKoS49WMNveVW/FKzLTLuW7PgiTsP0
APEU1HzRzy/H24OgMgH1UayDHn53ZtqPlYOiS1/Mnc3p9RLAkbRa2fmT+9bbU2lN
w1qvts8550OXfNvh35qRRmPcpz5AEtlHmzH6ud8yF/VYtBzEH1EY6fjfaS4KDX2B
amRMM/E8HSzY3kadCf56H5ys0aN2hE3XksPA5sNM3y7X+sG1aYFmxaUW6ByxpPhs
+u0Kh3sKCvUAA/8ttrjcNmsfVZDFXum2ZiAUervptbEvcBje+KvcXuaBB+NRcrET
AzwwgxJKNKuG8qIbOm8QiXCX+gmX7gNlBQeo9130Bi+j6tpMewudYGD4+j+MH8RH
bZLasN+jUusQm6xsXqsYtUrpD3n/Qq04z4x2NECgfRv68ByuY3gnUhi9uEfabUao
WllqEeKrrI63Vjq+8Zn926qF685Lmt2jfV9jMinWCh2+vjy/PxS9kmar0iM8ikEW
YQvx0ZymJfIr9zJ2OW2nubCZduXlQfiRjHX9QDVjPkyMdlg7vfeznECan/sEA5fx
UWUDW2e1GO6cqr/fDfnshp8kNyFyqvATtVj84wW0QXL1Mycd9hgKMyaNglrkZ77W
qPa+VOyQ0RcfafOVv2afjMGC0w6UNteoPT/Uq7P7KAKRyPHBWdmeyHc+OMTUhilZ
16Lnr2+LsauY/aycWhvR1l4eI2NFxDT9F+Nh54xYYOF9YgQJ5r3iVqju7RaNHfl9
2HRsYdfKgKMmHDUUwxMC+GLV0gPfwNw8bymVpDo6TiaE73a3Y+89i+m8R/3vs0XN
33GQxkStCA+HVNgt24P+WgHvIS0Rjsxlnw641JsonSLrFPsz4jhaHj+n94oX75hV
WMjcW8HlHt1B9oL4UvOolvNFjY1CRI90M7L+H+/AYcsUdZ/y3Fw6ZNiSNkRSPwaL
Iv+c9CylhomsTX53li4Cnp5dJjZPgtP3DCTLxWBDy5r2T43PHqxKAkndeOT/IiK6
o9/6ePnM2n0W01Vh/nB0ZKfm9q4/PPzN+XuslYGj6EpKJ7oqGlY3K3NniK1YhCuZ
hc7k3VtWjBvAULACrN0VuofQNzvYSK/DRhqK+uO8m1ubiOEbOHP+0ttn94mFatB2
sHDzxpdGbr/7mhIFD/z9PTKEYvIoIF5XK56YGAvqmkSlec9S7bRO7F4sSIgNeuAB
G9KDHf3DwsECSIq1Tbx6p53ZTueBN10cyBldPf1B7lhgjYO6w++OmGVhuvZd9dGf
TVzKa17oSyXygDfADQ+mb2SOP5gvxpg+aWdZIGTSKjll0xdoUVqa+D2y2M88Q+mp
X7Gkvd321zr+wMn2+6uD3GmuEnhWZ1eojNA0JJeL1trYgm356uxUoQIkp9Z0dwtQ
s9w3v4CE4/52/oRcxOpQKMOlYIsRLl6MlR1Rj3IIrLm8DphRMYsEleeLTtbIQ3rc
1BQ/dY+ubFuAOxxOBY+JpzAzKIh2gSidTTrkZUDHt+6+AVf8fEpQtIi+3nbHC6gD
Rn8Ltv3dxtqGrGLYAPsRF6p2P2Uvggkk1lr8B07cpzxp2mtEUT3jz0y7od00oBpi
WNI4v8Eq+26DA3TV11DHU3XRKIYVBqpnpmRq/1d3ExLLC16jOXbVzDjTWbajV/vw
hSiltA/qEqQ0Qa7XEyWgwcVmShhZ0Y0/JILr4L4DQZ0E/6XaA1WP2HcJm2HJlplV
2SG9m/d1NlZ8IwojdwIiM1ww5E458w84oNXfgtU8vECUX/puuXpr2od6fFJDPAnY
2amdQ0Za/SA6xtbwmQ4PbetxCCkOcmp+TpxnIVLWAxLbsztFSQps7xH9d+J3JqEb
8RIAp7IUp2x1hbG/34Wp/4w99hMp3Es1abz7yo9wAhGpJ45ktKQQ1jdD42hRj9Xl
wyR3K7bqtDqR/krx36a1ac01BKBTyYn648iMcoGv1Lqgb6Riqhc6eBaTcgZLNu/V
5Nw6boguE0eUakhZDppMfsxnElI4kGQiQYjCTU8s68WWFHeSOvs9gFIe0O2WZeTh
hHfWZ0x/KeCKwiOb6sGDlwRq3UqzrIXuoK/BB13464OKUkX+Pw3T57GoVy7oYp4q
uOqYHV9tgr7jswzJ4r2NYMG4/iP7Y97iGQpny+4pM1905nArRaQo9c/3yknVvQV+
152poPo4GWLoUt9IFUywMiFQBnjWQ5GR+E6OMkUymLgrP342SKtqWiLp2nmeLH0n
IE0eSmLkMunsNEoL3Nkw7KhTJGigSqX4RoysySJLi0k0RHcLK3hjhVj6kN0E+OAq
1aOvE7u8rMbhwxnFiGj29irWl98MKZ/mK+iaXuR6TMUY932lznbjkzL4h12dd62S
p5ZQBheQ24U2/mePfXWfWcdA7aMAEfPXVK1kwPGd3LvFT1Yo5QISkdLJGB09vsJA
/9c7NKmXYh9jOamqN5HUrDdo/DLU3fvES8jadM6isQGGmPlkIqW9U4zor3k6mUzi
caSeL4crLWUkywu+Uxx16rJrYUX69/TiSzQunmfxvfpxs+Au7GZ9Z6lOavkk0ssv
0sFc1lA9ABpTO7vPicUjrUesXrZwW+rK4GXGeKA/1Iew/hKay7gq9ffRDAVmXGj6
RXhCbuHcI7xukg2kw1XXwLC+8TXtcneWtdi1o4ZQs2MsksBYiE5XOo4QbxOU0vDg
3unh8yEnumgFGceuzX21JFXd6dOYXzgJ0XuOCUhJYFyvTrvAsukalHr1gGyyHATX
XAhoEa9czHPp4894qAQHQ9uTBD2YpRAyCKfW/+kKnS2/Djb20LvS9eXGnX2Rm/Cm
bfqC0wkbOXz2gXmUJOgu5VAgGdsU4EsnVAqiznIyRYzhUZ3tYxR7j1pUMgvCp1p1
bbB39rDlI8dum2Ab6QadgSdXSCDy8JlfXODWrhTgJQ9HEA0cO/5+eNdnyCGSKJkb
q4o/q5HJIDzmzxBqP6Tlg1M2tRg7ljqIjEA2P9J2Z+Yr/GvzIylrdTrah1CP/N8f
RmanO2o/PG9/hHFGnFwoc6r0yukLRmwboyc37DL/KQtA7/y+tLUD6bw4/57d/UBy
1IuiJoHCnUgef8CNHjaBbpNG6VwlfWfpvqSSKs94OFDAscScFbeFFTdelTw2GQqS
SIK5Rw3HhlJFhQS/rbVeP9IEfGbfXY7kJIAj7wstQQADmQqddJf3aoYCuRoSR5QY
rVs9QxQCWnbEqR4Zv84iIVIZfrZaYFCvAbiBsea37VQJnXCc37ktcUBoKqojHsIM
0FSooRqk+igF8PI6/re4YeWfSPZbR6QBuIQ9Zn2o/2Br12zp6odioZwzZJzTWjbw
hfmPMbbJ3Cd2/6QeukfMd2vVyC8f06PWMyMf+oP1DIFCRj6Nl0iYBhRyNjwxsRbR
cOIwMU0X52IZ0fLhXGF/oUs1n65Yay2e5j56DUGKn/w/K+C9KyKmlEUN5+otIe1Y
spbKWv4E9fY2KTTqsgMb++CEPaX1Ezu6pJH5ana7UT9k1dJZDax/vUOsjWG6Xn27
LtDS8EpNpdW6siDh1x4TG+agUiIXgQp4rupyi1XOe2OymM/SFPl3GUEjw7QAMoPR
hQOKTx5ytqOL0JAi2pq5pTg+BWDfD3MCXYx7KnNqlRFckPYuiJrnEzzX+fu73T/R
/F0jQAQZ/vAdKNC+pradO8r1yv3vyPpwvtPVWdxJjg/7yQ2hA4hp+Ve4dkEoID0F
nNFMbI7ciXZYDtk67Mo6X8fXI3CQbTi1wPYDFb0HU4Gt074ZqLf+mkcrYtniYT+X
TMDGEb+VJMAa14CqJSv08tCKHqBk81HoLs/qHyxV9uqlpkttz1RaI8/Ubhj7KwR5
xuoEAZJxx5MYL3Rf57udG3pF7rXZ/yqAhFL+4hr5reh20iGUbJz114KaFCkMoOFZ
3NWzcZizOoPqXx3DP4/3/Rl4NN9/VoVl9UFp5sJ/3ESNuql9DxH8k6ffLUoQ5D25
oro9kqp9l3EbZCpOknJVu7USzwTqgNMrBRoXkxe/2BMuW9ls/A7LJdqJeIvApGvr
lEjaEz/ROfgJ1sHgtvQvQtOi4PBmvPy7zc/Ha/XWXQRvWOergnzXr2WJqAnlb+R2
FK0ZglB2/vamFUKFpUNjL8SUA7AU2loGj6TLMY9s464sKh2gyCtyR3FBD786Ph/z
ejIy+JTEvlwvG83d3FU51+kit4KL0LeB7A6QUM5+MQ33iPLQwTJTayZha4TvE4T6
NZew4iYHiHZLWUwxr8hKVZHIo18tBomOUeVOgOjhS4AtWmdXCzwaYxzXXCFy0Pcj
bUXJ/Nt5xTHzRy1YXfVwMAZrJoAxR9BFV+MX1uGUNKPnPn2HR4zAWIQcZ4DdGMEQ
WbuWi1iHpqLq/f849yFzEcmbDxW0JeC+ih/T28dsWjdP8c/kBj7fYlBLtmXzZRfB
FixTYV6NfyrM9MMyajn5yEg+pwHj0lZQ+Sw4s8FkX/n0RELG/5j1kNMgI5iZIYVi
+gQh+a1IItH+FXRm9dNxDTc0eLGCfN69E4RBCN+fVLx8K3e0H0X7QJxyo4e77YEy
ZXYgKPoIvQN5bc/8rx/sTa3GB4relgWQd2q1FEvBsiZbCbxA1ysTOM6ZBabmXK5d
Kcf8vdJZC7WZOwU3gjb2bfl2zv18OupjKKHTuZdJ4O8TBrZoLRWE/GMwVoRCOKex
umbBAzU1bTFRKfQDct4JjvO1oo2J3BCWsWy+y4BIsA1krrk9cMQKSS3MHSP2d1FW
QkfdkDlyU749GaLE4FTsqw0D7PJhXttHnbDfHSxmamQGI4iO0qXxTFGtJbFVEgq2
k472NIHjLTB/TUggt7RFxmF8eZn359fjaPaHczaRFgJnh6lVIIHQvGHqKwtFyvcF
rWR14+uJR2K1rjZD5afnW3SjJ6JkMF7dedXsvKAFMMRFUXhcg326qGJCj83sEoff
VYS644HXdwemyNQvgNGjDnxd/64wGZ1KWVSoKKDNfCxw2RVEW9MN82h2daYndzwo
aCwU/HrrZ6ug0i+fdwFUixCcaw7ee5TU3D6cKgdQbjio85MUsp1hKCWtAFa6qPat
yxBJ3jZ2SLS6f9VoDv45kUw8nuaO7KDOtKrd+ipbwKKFh0c/RRVomSp8/qUJcOO2
jLd2lGB9WA1/85gjutRIZM06mmPVUDv7PpN9KalnW1JBNZFC2yLjbSY1AvNOup4u
a0KZQzP8/VzPWIUBDkNUaJXgIxC4aQdbEgS0rXFuouPq/iaZB/+DS3M1XRdwz84j
ujR7icwOY7Vzw9tOx2Js5nfmx2ZlVyabQvN9C/o5nCixSGNvfxrYQccLkJveIfAT
Q3/xtv0jdKRfGrENnTi4T6GJ0zwc2keTzRFKidRA2E9WOZBRubrW2nKYeENqEevC
my04685uAeybeTcyTDfnDnTkSXL8PFKo6DYCaZJnGVczXWQd9edXc0DwyRYHbLUy
doTXr3+Dm9RN0B8A4UVXOfHIiLycp93+B05TJVVy8iVIj36CZs4MY7utK28XvkXp
5UggBCh3mcZXhkNJ5zg0zzphYVXe/eN+9D4W4RdyaqDaw4ABe7LbN+/jCzlg7/ww
Poqnxor3wS7CxVY4Ju/DEMgIkJvWNIE/LY82uRHX8rK3accnlE2ZJ4eZ9y4jOkea
k2NzMIIcmgrvnNLGfn00xv26lvw/VD744fFmOVilBYan+8QKIdWijPcrHxJakBiV
AYZN1eLeaVuR7TxzsHxFUJ6uumCEuINUPGR2Yi95U/BzTf3788Y7Zaf+irDkk37I
C0RFnFFMHdxb+Y90TfxneWhHRGNIQ0h5j8cOgIMjRV/ZBk2yKhTP+twQkO0nhRNn
36q/7ewNp3WSQIqd9sxM5EKR5290tq+RxIbSLeYbOHYRjdsnPcAgrrZJKSklcC50
GVBPvWZ6X+hNJPxCWFBYa/vFycGF/YjLrmzLlwRzibeAeEnubQ+KP1XjUn+TNT8m
+gwemV9N2oUw370gmG252bvxJZSYi/fg1caiGOG8Ah4w26kcjj1HvHjOJCN3Iupz
Q8Pi3TLgcj4iUXO+XO0MA2HEveaIfIcnxHzSUBDKIH4sG3HoO2wzE6HTcnIL+LR2
Bs/y5ds2CLASJsg/GTjijZEI2+yGNnOe5XJpnNPEgti+g+vi7c0z+nUtEGWdZfZL
tx19gkLcx/Jy0145eaOo9iGdRX2CfMPPfRGysL4J5QI4onnlHMpzNwew8PASzWWY
7PmgvUIZPtCgFvEW6J1NR6ypD4ucS7JBd24O/vQ7NY5QKWtKqRwN719Zl9gx6WQF
sh0c01qf8qAflR49j34dnm6peB5MXS5qkH4qb32/E2cXMVLbBMYZdBhA7e59OFtV
R7kq11Gu0GC+g20pumP263w0kSmaZDOiHPS9pdR3/+COKxjYt9gWRjxtjCOjg9zQ
ufYTVh7WT+qB/zjN0kQOQzSoquM96ksbhTHuxHZcP4Zh3GLldHmsDhpFOgWSJN7N
ksDOLF42uawCxhwxp1+Cf4+6H6AMaPrd89IPfXqMMP+VFYj2UvXQZtTihA5zaJf4
zbJkQUgcL9ntXEkUGo33mlH/QrKWQ9K1//RJito0hYXmczsa5YeXkESfIBxTMXva
qchYdmIlAMev9NDIArGOAV2ME01XO5eYWX25FdkTQQgX/ZHJ666AZqAklXaO3gTY
J1yL0TLeH8sP54ZI6RG/ga9ZNxryWAsNwD7YIXCCOsabuOGjDUetHDEUgme0kWoe
akoT+eK6xeKiu6v7ovLMFU2oaNPOq8nUcrJdBQXSbOzAWzszvdIVXdAqKYJ1b6x3
Sfj06as8v6R21oUjQOm75axbZNgfmPXHPgPjyO0g8d+4vauVWiippWIiwcla5lJR
CLr5K1sv3imhSHfDu0rXg5FeaHUJ1AIWhg+B9ZuJsq+iIgm+8ww4qxYOGITMH0tN
aSnMMRE4eM7vk/Dh+VqRwqgDo+rLiJ8xmHWWg3BCSXZen48ZJK4rpR7bWGKHAHYx
tOM07ds1Ie6SV4QjSBnXZ7jgTgyO2G7238lkr0/AHzZTUMc2gI3dPdhwZ/XX34dC
ZSsW/Y8uEfCEgBYIn/NkVqf8pTexqSSLl6lOcagHRLrVuWJlCCxKUcJFfvLQYO/P
CfxSSoDp3xunZcyXOiyajQYBZYC9BcTjdZx7m17eP43uNKwbus7RSjtKlTpkDfTm
Q0EbPQ59G2X3xR3Gc6NmidGYiCHZJiYl9uuy7LTNTk6+lUyOljJpwQbDE2rUcMsf
dCeMQ6yjDnzLbUFDEmkl/sCR0Pjyt/mKk962UDKvslSsSZ2WV1YFQ3vY6iVXDkeh
0plD6I90a/E46L7VnLC6Z+hydWhB5u6t70uEkPYt1sUjSGu/7cx5t10nnju/Hq+h
YMkG/CWt6gsgKkPk5T90WvIypo9GBdaAtYRv5NSiKdJRx9Sk21HzKmJjU2lRxoCB
mcnHLbPfFTMqR5HHhbEYo9zsqLarAUnAVq2aVPGf8F1Hl453OxeUS6u3Rdohqw/c
gr044HlMB0frygrlk7/X7w667NU5fB8wWFjj9mIBTdCOgClsGKV3L5QV07T56+k+
vAG8A44WNKWfdNYtq6sX7AGfhOKMUs8MG38UlxFsfmH/BFu4LQggYkkcukMt6E6g
KAQHpktLbqOWUqpAyeCmtHTEUSU3ICYsEMNZH0ho1/4QcqDk3v7WJ1hTHw3xEaca
idMhD8fjO55+0kNp7Zl5xvwFC6xJ+LdmpwNF4a4f0UGAJtwqOuJ6lATlEDMlYy5x
23snqsIaGoXhBla5cq1Lzi7qL9pVZt/gWKeGbY57sdNRLjZVIhWsEISi3pxxMw7w
8ad3pvDbheN7h18AOECeiU6FJELMAzsXe7/Dq/PN8maywYxP+cxac46lWwMs5JII
HtOR40dtyhFT24UtSpPbMaL50qIR3ul4r+nYIk3TYxsQsDA6K7z4Xdh1UEHXXJVZ
/7/WdW1qn4tdCuessz93jxS0YnOyq6RZMHDTGjfMsBDb8tM8huVn2KZq8lGo0sZm
Vt0TiqSCU1+Jg9Tm7vaO1XO5FE7QPxNG7JWkSdDnkXCVq6+e8anAsYMg89ENnE/o
JjgSdfBY3KHgzhKmrUkkgO6V0SstgQ71j28kvKooMNgOEbZBIr5Kw3KclAc+SYKE
CKTA+Jhkmapd2g2pYd6puSqFub5nQrqzavs55KfWLxgdTJLr1hC+GMqt8mKbYuD2
SixzcY1kSBt+gnbDwvp4mIyd1t2sdWtdFUxu0VrvU4OhxGSRLGZ7Sic2IV91/XUw
EQ8Shen9fsJDoom2b9ekil0IFEBVn9ny9//6gM7HyJGwI5G8ruSOYsLgSQP5ByF5
zsPsvjoUC+ImI8g5NARbLZ/s4pRfyd4cwWAU3dSh/zO5Xm70txO69BksGkUli2n1
3+WYzl7VglVSkkQ27mJJIwcD7OAYlbt6rzwKxnNO+EGqCu9xFQ8XpuuI3O9bO3/0
1EgQ4q9An6HQ0BW0t8nfK0Kzeoudjdka8fEgMr+iqdjcIjXYH22CdFpotuV71ogo
ZdCsbpTjzfZ3q7fRurPiWeiAXskaHqFcmKv3gLXPkKySp2YDmQ0lXOs+XvDC9iOw
ERQm1plmeG20SqMP6Fvcyly1OO2jz9uR5q7ItQM2FfO/7/OHGmuxS62CDBB3VdLS
Y+z1TrDW7LDWymXDMOBn3r7oOSoo+T7QQvoPyhTIhJLh7go/tsLZoUTE78ei/Wnd
UmIFbpVHMtsKgM8Q/taR6fik7hM5rWcObwZVgyuOVKqJ230MT3Y5toIAZmPlPDlB
Fr/zfxSgMpz/k/F9NzXwnL5N7mbYq1i8A38mrt/+fvfLeqRivoBiflcDboJtr8o5
v4jRnGHe9jDP2yZEGh5F0fGIJCfbNRc/PP1eO8kwirq5FCT/7AJicy8TESHJ1nRA
MT5uGMRTUFc3vZoONM8qrDg4CiUAYbJrp5wUUSKQzluGNJab/NgmS+2S8AU4wpzU
ryqdGZBLElkupHXGddG6vZ5B9fqT/U9F4iuJtMfkWj2wpktJRUFCI4L9Jd7nuB0D
pJ31ny8KjHr4zlk2lnyyqHQsP4Xe00TZQCFS9BTDQc1hUIGN2nbIK2HjhupL8Q7Q
YYRubwuTM5e+7r2vYc6mz5+AqUmDahhqTKGBMnpjcoUbBPYEf2qWlJATDBcU1VpU
mS6ITq2ynst0iiTLhXM/zD9HpjHaS3xgeP7TJjBhh+An+bqk5uDRWXK59YdlK/EQ
48zOYXLj0JQTlSLKxbLzyDfCVE3m7nzzrCD0Ksrb2cGIqNGDGaYQznehXY0wwx6P
nIDYoUR/ouCgD19nRoT1ys5BhQIE/oWlzVrNDA79XcLk4+QjRn0RdFRtBfN67nGr
jQ7ACXOv417btaEpWBTTTRKVPtYNLNFBLqz2xg4X0LBryt2oVFnAa4T4Da6xZ16a
vkC0gPEYWiriHeqnfNaakYw45AxQAN2JlehZM8P1GTzVzJ59aJlloFgziyMGUAzS
wjx1tRjX1dpYp4UqJ0ynI0vF1sOXDSz1tkwSkmtQwG4Vvr9T/Wa73XqfBnxVrBTC
bpdNCLzxL8by7/ukuZ7mAu7putabtfD8nY6t6WlbZP/jR1HqL9R5iTaCMSSzblx5
4QRo/+g94zHGoehmgIUhbl5THr/JGq9BM7fGOJtmr9eHix7yPTLSF5m9djRQ8G+i
y3ZE2D0tOVqffimYJbDFfFq3nxGNdFxzvOtZFJE3c1fzE+5xU5WJNbcNnuMTz8iK
QQ+sPu+cshyL/Oy2+dm4akfB1gVrnawb6Piu584a1FMLi2hvGWIXpFE/ydFaKhIl
RLfLOocXIJ8pFrFp5kRQzolrh2itD29LVfbADYBzIJmOyCOMgKqa3Li/f6BwLCRz
fkPxfJ3F2BnO0sA5/yd6VC5Qplizbse8HsmKRhjUH2+tEnhFiQ1lQgEokcdHBFx+
W0ekyq7Dr44TiwfMtD0a0BJGK09ICAGOipMWvNMjpeSL7thSN5/6jlvKKysi7+oo
OlABSdBQP5imxD3N0TpzjamHDILGT89TvuKoiv+H44WH//uP4wubvK1KhBR3ROGx
dVYjaPAxSlXUMgy1Al/aypPb+OIrBggaAfWak9iCx/dhKmsmuClav+tT+MBTUiE8
Qwai6jeSLxzoSh6yBVikka1LHtv/F6i8VWSbRWWf1jpJDO27boxEywmf9QRQah0X
WRBKJyvPIvLLpeQE4GmB5uTnkpnvzEtPJUyRDCui1NWtXb9GLUSQB0NUURirA67m
o49e67xCm+klYoBR9pVgub1YRdk2wBKLv022NB1aPyN8a8rPBO3S5TRlUh7HyeZr
LQy4/3MbwGQJlgJOcxNwdGkOCsARTPDdTC3C67F+haTbs/rh868v+cK9j/okvCqR
yyVpGWl+OjUJh4l7jexgZbpjxPwX0aGevJEbyrBhlSwBInfeYDl75o/ck7TA/EWC
flYxyPe0NdE81OSI+LKFPTYjs5WCDndVe6Bc8pE0+s1hpYqiNoVu/jWr3uLMZqj8
FwBK4bz7w16nhhWx9CY5yF5q0hwkEHXNTj3dH4y7l10dHGajehI9bVHwxRbf3uiO
S9065engN0BNQNWeQTjZ/efl2TuJmymD7+Yps+6H/fjdOPAkyywsJtudN6FTtW2y
Uv92IcemuUAtoPumAP7n+kfhbOhtkQqY5LnAYv1JKlB4kh9AA/VZK6WemMut7sG5
mCyKalSz7yp27zd1ZNqOT7qPsc3IQCHqY084EMuu4k9jVhVBpzPi0M7iFQ5hlVVp
qZKu9kLzpkpda0AZbOPKA3ms3hsjS12I/agWZiN+knJtxdv1Sq84zGx7Z8tcRCfL
pL8V0J6qypj5ilVnTWj1tXb9su6OpM80ftdxvIb4RvKIdWM4dSLAZOeIOJr/aT+k
a4sbRHgRTlWXqEVEAZCZUR3/gh9RT80meWcunS4oMarCNhXFlIVNY4P88Sf0MPp6
YgOng+353Q3iRr2ltleHqybT6kLliMWuMEYpu9YyFoTBJmf7AGkU2Tg9nVXQ97iI
DLqsTaAiXnsNjGd7koaQDzIc38QBtHne6DpoBr92Dwqdx/yveZveGtKoUR736RoA
pqqsynqITBu0zvdbkFhmR6YE+Pc4ZNSyELqgkiS9L1OmKxPNMtbl4hjdn6NGnF5Q
VG8y0OsGrHkzhZ8Wz6RZa+2QM6+zjeg/hYXPnSf1Ql+9ZpQTaECfkhRDAH1PdPED
oxlDK1STTukX+M17Fv/eD84+fkVJGQiYnJZwULUK+734ywOOtlfeF9ePZ7O3PGTB
igGaI07XE4Wgo/DU/4RpCRrpR/j48kZyLTih9B+aS3C63nbiSWrKJ1TSjCX/c9HQ
mh7rNOJeHGIV+y0f8HieezTyrUk5ShhbmUBgeKXXbztnZcixSO8N0LiyPTt2JX8M
McL+tDch8o7P5Mn/ywR6XccUmTJubKNixrYmyPHt9GyqB47unoL+DVPD0evIK4ql
0AoY4nZBvgYtTm/QZtcMEgKCjTXmwfMot9BsCenQG7u8g+u1ht/MofZ8zA8t6Q3w
NzX3KjI8X2HaPu3Ex5B4D+o2cz69kttqjQVOBBN4nqCpte/UTGs/cKXu3vm5ejru
n1pDO8+/h/mHWHrPU6XtJmdBaNeWky0zAqe0VIDCC6z8YDEBzPHwaHXm9/pegMEw
UizFdAD3gVSaGxhTy5MFrTkR2XCeH6wkScgPIo+O+rCguJ2BIVESUeQuHZ/Hj4gj
REHpJEnsDJ41AuouC3ZuD8o0Dsx7zR9IxoBYwo7fVy1DbMiS9iOEI4WwjIujfWoj
RBWcVMtk1jXz4Pc+ZA/TfPht9OJ42QuLlx2xDauAYRYpMU3YB68aKJzC0vow8aUE
FYIKYrjpDZJ0+eHjYCeLxn0769KgVeT7hZfxFsu53HY8Ymans3nwJiG6aUEzoKN5
/wJQAEA+1RIiKGuAwyNhUsI/tdEzOfYPWxQ8POechMWHtBeLVbZYJ9OKRAYgdM3y
GT5NbLhkXd0aUJ4dcTZUDS/ftuxSU0gBVFVpcR4v+Rm88cPB9z5eQvLyKs1yPWuH
gHfVzIs6rSyng7P4dCXpqTxTFB8lAaFjoPfU4DtX8o6PV1KbP70SZAvxDM6hCjHq
yMHVcOFOUC7hbWMbxd4tp16h5GJYUiVXxmFtIPRoSVEX3AcU83+OXE8YRQR5Qo5H
H78Mtkyd4flImbEndNx9810ZH45mxfYwO1xc512av1uiHtRSVuMma/nBjAwMWONU
pdma9UEfFov/ykw9/6Kv0gnd4eOvrvOqu/CxFjOX5OP4Xu1GnTVaR9DJbIGc+7Tp
GXrLnpxEFxGtwTdNDdEcsdUxhTJhQ7zXWGX2GNx13BVmjW+YOS13lFAz1yYzgiEK
i0uCLloz8lRy/EPKz66bvwQXP2JBHLoVXc4ok8Qj/Og+84WQeYKPQR9ylysKzSTu
eJnpSiS3aHcPxFjKuG1+NJZLHPqG3cLB6SyeDQ4U9XaI4nvUsGl4m2g1iUUlF68S
ecHMpFp2TxOJleXhu3yCX6nqgCiujzP5YuXWE59zCDNx1mWlwOiH1FU5nTs5rMIh
Dn2+8UGyt0YXGicwuli4b8RXGbFjBKdfHvAvHLHyhPm7EUrA0on/hhpNrkfigZYp
mvmnI3ybGS5/j9kimWsomT+H1BVAPlRcr9yDyNcQyjVcnIklDPyRk8fTX1nuDKO6
TbaGPwhGfV3GFpD6HnOZS/VHVUfsGGM4Q32QE/tYNzboiMWJcfA9ycYtC0aZKGUM
zj9Q2qK0IlFBsSoNYOXcV7ARwgXiXBTNOg+xFIRW//9LKCXOArY7Pa2hgpzkwkaW
r5UervO9xWcsxkixjsjDxmN/p8GHmP+VeNB580iRDFBq80lSrcmQltHVummRnHLO
7cyPKxcd3KIdByQJaoLYpy5kmIWscehjFZLnFWJEgnoC1VtWVyNul+Ewogs4bHqv
GkrJZdEI/I2r4DWo9WoMoJ4JXr4TSOE4Yry8bM5PZYb3ldKYwW7YU6BU6K3H6rXR
x0fmFZf/Vtw+cBCrtPO+k1g4AO+7Lnmw4uF/3SKD5piEo7QVaEsMb1hiusWUV5uv
HDx+0f0ROVZhO/KFpka6sgtMbgdkphjmJvR8QsXXI3XUgnL/egIcGeAiNLep1HBg
zeydHtfDoPec8jkNxRhbi2ZnAj/Jdm6CjglAMe2QroMnyg946L3ZSykj9rm/wIqK
oL94TdxxI4TiJeBr/JN7AshZVGP/bIJlGHmf/AcCGnHkyd6BzlOjUEDDlrNRX+z0
6h5uzxmvPUcSBeU/lJQYfMdn4wZFkDST2hDlT5Q2tE/T03kq0x7P5BgHeuHTK82Y
DNaqv/Ug/SLIVfyffU4rS8Q3/zX/D0z956N4ILLNQRUedofNPQaIjDPghHepp8KA
E+b3vyTgJ2zJrO6WnrQsAaasetZDV52Gd+oCNfrX8NoMF74CCswRdbp3S3ySrzBN
jkzuu1XvZnMdr4uL6Q0172uUI217l2ZTjLAInc63ezOf34cEBqfC9UxaMo1Xg05C
de0Rm9M3GL62W5LpXVLbsNaC8mUagjEL3ahtoMUFJKdiQCedTHV+Z/83A4lfms8r
2q3k0SZM7S0VbwRVFyYzWhUbbCYDSiA1M3NLiT8yQezVSZYaGypLfDASL07Cx72x
ymCq40bahc/PApDTnz5RTQ8I4qPE3uu8cBsFnfOOcLOo78b9yGqabRcx5XstG1dV
rxiNpZvhqh6HyGjlb+wP1PazMKx88nQ9QIW2BsH7tWnV8BB5XBXscVPHzzM6PZD9
3faA8e6TLXTyDkeGSfiIdkzb2GClet8mx9UjircnSyPZ0b0S79/V8QFX/JS4tLJ1
U1DTlr1kLWuMixXlnZrOYsCCTqh+knyBQvWwARn3udmOx+z8LLHkFrRShtlimnQR
NTfhAyA2tsvZw/rX62FEPxCcxNnMN5oaOANSu+Km0u09rXIOGu47woXxr4LrL2If
HzsxKLpAW9ldFtRhPWXXo/SK05isZ4yExfgCQ3EaqC5J3r4eubJrlpkOdKy4XMaL
U8nf9QheB1NRmgtDlH4oG0YJRmR7KihG7pIqAANqjht6uM1JW1er6ZTo+aZ3CCUd
IWnkEaWuHt7Hpw4eDdVmE34YUJbmqaMBGT2Rt/YMm+hPPuDmuN6XxDY9NhgWKwIj
LCxCXb9GEA/2lhLH7hpJyx9q7mBriAoFBacWeuiFORu6+0ztxWNsdOqu1JDNfIg+
3VNQMpDk1fs0NKP8CE4Cz7xQZP+KiAVX6AOwM9kOb7Lv+rlX8oYhsdRzJlC1XwYe
qRAu6i5aGEebB0sNNVSj2z7XBffDfPyofSr10BVVol7U4NQwCApsMWlawbG0Xl03
zu1V3kZkS+32pO3jqo4MgloHGoizWL56Crnpwvk80OS/gH3APLRLB9rdCBkDt61R
woUtiOCPvPi+zak99Dr/e59fiK2nPuqXPzcjgoL9S2WvZuxeZH5NPSDa7MpjikDL
k2WpMwbUtMpISHLYjhKGhSDFPWqvhDqR+oHzWldVmW3RsZ24eRuXbFEHNQIfHt86
httoDZIa6jyLRbL6njLN+QqHCNQE8CXSzp3LWKGlPQnV8xgevQlQFWD+WzdBiwpY
I0nBT8KFrK/Sqyfo+jjd6FyCVGngOwkVdNUFlKCQaZ+OQOePvtrfHav+FvakbhnG
v8rKU05H6dOkGlMfqVsrQUOITrc2hf2ZNv1cvS42JnauVXiijgjbee2dM+GyWrjM
Tnb3iKiwUNW3kgvnarz5CZHEilFuXTRPkPAQ+HwWA+sJzr4jtvEaKAC4Pms6PTew
dTnOCCrpz2+NMdHOkQ8kcJlLohOY1PlrqNB2lNMJ9rEU0pJpAykf/JeUkCoo/QJo
s5zo8xnyFByZKvHCpE2zeTA0x2fdKKeS0xHpxGy8daP5RGLNvL8VVfzYVX6JE41v
XGcfHDD9pQneC9pHaD9iPkLAwNGHUKmWdbgaeDhio+NV6JL1PHcSCOv0On3KPvkc
vVSuD/3rRXxwvdvrFCkzZMTkvxO+GeIU1S4+48oTT9Cr7IUT+iF0ffDIvkN3UipW
xVGvH2CB5vP3tERJ4MVbVIuZArv1+S1YyJh6mAphvPmK/RR3v1Q4YcuiGoRc5BJ7
wjcGxARl+M/Yef/JwR9/pGnSYK5yWl7/mFxePKamaujMEHdoCQXEo1iwxTVVQviR
aZtjP7ZLah7sCrDzncf+iAGm6bGkJ/DkdB9nfuO0Te4nnOILM3z3Uk/otxMWWl3/
TFuVruoNFJ071BZ/KWz24CB86oq8kxZcKW0X4piVRefwPXonP5+Q/u2AwYHLjQpJ
25UmW9XVcH5yJBYDJtklVMDkfgOJdNYzbFAD58Vlx3rH0+mCptk7DpO8s1+3hJfd
3A0waiWRosyYRI1K0/AaqVXPfYYn6t7JMEwqscIvfEz6afnoO60NzTFJsH4SfaSi
7hn7H+Z8+ULz7lTXMPQRDB+BS9zb/OPflaGvi10VTXuvBvUojeouLDOf/FepGiJJ
JvkkDT1gZsDFoUf1CIGJRLeQyOfWXyQaP/oABqEF9fAY6kKcuNqdKgb8bVwnv67C
Stuzu2/MB1p8YMbmRiyzCjg/LSrhZpAW1i106wD/hIiwHKnienUEjbqvdCA/OPZW
O0KZu7L1cpD+JSPD0fJ1hPvCiGOhqmFwyQ69rc8anAHy7MN7grlk62+tWbW/ANWO
h9Um8d6pc1Y02R+5DwHZJ9dHWYy30bCiIeVFLLIxEYXBMNYamzTuLY+7Y2smBV4A
uZkV8b5pzwsyKG80gcS/i6eFThVe+YrbTPevP5ZSUxVFdR24AhKDH5D6+38V8yco
mYIxYaQNfpSvi+0dE/9AazLa6jaR9T+R8ADZ4nB8ARXvTRzgkTW8c+Vjd0pVFDW/
4g5W5JcGJZaP3vVaMLEn0Cl3tT2XMsNl1eT3c6YirrT7RYudC/dY3nauCzABGehq
ijb4lr2zoCHP/xXVhfaNkSccfqW+9gJFyvlOiuWW5hVgPIkDlGnSLivKun7uwDZ5
A4I5ghmOJKUxm54GuaR5CVcRFqE9woSgPZuZi+I3kXpYK9eY6aHEYsQTV4PTgNHY
+ozrCkYseNPcmT9OUNBJK8jx8QTS+coMiVgbP6CQ8yf3zExTeUU+TA4ZfCeUy2wn
0n12Ll3EOF9NrA/IgNrhW14NEVx2KKJfhaKcs4waUX17hNrayp/Z6n2gWlx57QUY
eHHMOgjWlF7J/fzpfqe0RT+Y6yY8XRHRIy3261vUt7L4z5BqYvPHw0fRl+Z5FqwA
lu/XTnzv1HjQ25nxHC2EORvKnX4JrdFP2dPdiprxUnr8BxfGK7OCUCD2PjUP9AbL
y6TbKOgw2CDLgHtfQx7q4nzjpd9Wx7YBFZDsiBE9SItpjhp5yPkSTEnjSAkml6bY
BBeoywi+rb8V+tC5GkWpTyqIRyHg6L2L7keA+ErwxsaexDgT6yRKIcgXlWmXBVBj
KfX33MDLtJ1byUJ1LjveoAJTe/X57yKBGsvSbMMkVNSjhiQSerbL9eLKnAG3jh7h
qxD+JIypUTiPC0PTSqTdt3BLdBHz8ZPxeu7NnB1J0HjQtuMZjmUuz8AErxNf5sf2
yUgMINahBoxfpmpk4FeTwQEYueX+kLWgYyd6oZw3JMHw0kGP8jv0M11Le+HIyNSf
aGDRHVPBLFs4ntvU2S8unWNcxyCSA+GZLFqetYo7YsAOMWjwegvXtHkSmlXoXapa
vNls8CrhhXmN0Bvg7EWeNCxtc2+UemSyFhsRcxxZJPcN/knRUGmWY8TYrybpi8ww
HaCAeuYFQZSiOcyE6tkIiAHRF6RsBZik+Qb8DGcaX4Ag1hTVG9/2v735ZIxnnHIv
9k6xy0cJEEmtOO2/sS9X3gPY223pfiCTY42acJZcyiVJyrxON2UP+bXf4WZOX5Hm
xl9WwczTDXZ94yoPKjSWVg5D836arXBvksexU/Rgf+taq1aUzfYixNChTAHLsMxC
1J2nrOh0fZ5CYcKTH72rnL81MdZWC0dVyYP6N24x+QKWj4fvIUWOCrqxKFj/ew3p
jfK31cdhoyBXiY1zi56rSeoE8d/t9Ds1bNblx6R3RTJ11zIG0TRcPszdT0Ri1/Yn
DjdfCIEu75wOi6bf6HNRQjAfEfpwLpKDCZpsUvJglTVq3IvwhZFWcLDd8Og9kN8D
8+0uAcD8qtYwAZxW4a6WzKFJNkUhCfQMDJsLcF4YJNfqyMrOb0SUxdeLzlQn+Ahs
DDPnWmm60+uAkTsRupBIYTjlm/D9ZO0AJX2nPRzB2SNw5zlj9WBSGkcFoPOgORnm
OGctp2rUY25wAUL9PQ3u7G20n59TlHqsGFVP2Zo7eAmXe010BtikYyvDWpf+Tzzy
1xAG4id1bszRjv6kn0RjZXTjZFK/H75uuG7XYTPkZgSjnJ11wbSvYc/CuLaaUQfZ
gUromzqu8j6po16Jp9z1sASwdWfA1ZcYaeeCgey8jZBv70fy39dtG2ogCO9wmQdX
9MWxd5yh8jL8P3EgG5lEflYvA4nNSKsW1om+syB1xqouTnqII0wKHYNvYUaXUFdD
CKBvLtg+c7h52+S8QPC02YQADl9GPx/UHDxDWfNQjUi9FpPAXwJlC07iUGu9fIaf
W1Bu8AM9XUfRbQ7WiA+GrUvU23FX1H1e6zeolE6LhnA8BLPBzKF+UepLjlPJSNM2
Re7YUhEuntcz5xbneLCoI84T2wVy/3zSoPDV97GeLvd3NzDRLYicb8aMlbbWXZAj
KUs1Bp9pW9gOP1a++ZVKVnI5r5lpdjClmGdwfkxqQpRczg/km5YfghQ91d5ZhF/3
m+/KRkHuPShXarE30PaKE8Z1vYvP/68Iu+gIt8mjv7YuptdtpTNXuO4NxzLfXLSq
Sb/OiSlNEMfamcKIespqN7bzCGpF4nYO+lYvnP3WD14aSsIn+ggRamC6Cv/oLYDQ
pV7seTD3qs+FzSREfq5Xl7q8RcMPTdM+udZYOAyrX86vwDiNu0XWCOcMxGE+wank
tXUP4gpgeAQEvAGn+D4i9F6vxyjhLGR7GYZdZYx30ab5BaQL2fA+1s+0NIY17CMo
bkdmCCnMy8DS7qGHepRZXfQBFp3oLaJqkELz1yq2cNa2NR+5Hb+mBTdY+88SQElz
iRjTQk15JLkTC4Hs0Za3Yzv1ac0oVJlisOtlQOthOqk2vSNF9OztFeCi2Dt/noW4
NvUjGOzH0whfS941RtM0UNDe0kdCfcEBdVhKGhpc3ZwaZXx0rOhVGjtqN7PGglls
9Dgbj/afa9Y1tGp82uy7uI2FD9E1ZehgHI+fXLChxzmA3WxObbCJFKO9i5o6rHn6
2VCFKHqWhjK1nOGfOseOzctFagINQXVASLc+KPUwLqQgCWK/fbtkyvql0D2folMt
RmKuLbJP5SV1wDvrL/0jR4b5gVwybqzp1pfdakt1HvnpYgQIHBs+wDLwoWI8n/yz
PEInMK50B3FIVnaUSdCyJmBR9H9o/mSGKkdfhmZ0in442bKz+sTmqw+LqWP8i/eX
iznkhT46H7slsf5/ttnR5gSzG+FPLQVm7uWnTP68ho+HIhG84OLNKwgtvdkdq1sx
dHAe7muX7ye9GUtivLWW4S8MyTafrqTP1vWuHIZ66HSXfDIbnhFwus+XH6ehsAS0
5GhP9bXcBDGHV946V7oKmMFbzAJipHstb6kvW5wo2+OsaawxaI9GaWviQUuaipTl
TnhRQGeoC12jtRnZL1xFLM1riKPl3RLCJOo/x+CfN+G1F7BQKf+qfBbfiDJ2ArCt
LKNWhVwq3V+15LtwFKI+T2eetD9K2/W8nCzBmsyMRiK895IEm5ieDuIjgWdW/6sy
8HKCSMYj1ARhsdtsJLTrcvE6QlKKhOixBTocoHPQ9zGKS8KqCzm3LJLPAU3TIDoC
W8S3nf+ermG9QQd6NpgvDYWhU9pDuyuUXz/DiwtPhqlrsA44FPuMEFh41U99Qjm9
kVP7K1/om0s9aqsSPIAto+wCiBN/cRc/QPj9HXmsNRxmFpTcm2Or4/1OJwl3eiNt
Wu28r4VTE1pWpuMtsdaXF6kY65LfVpRmHf32mh0JXlj8inn4nSqa3vSB1+VsiEsT
RT6PMtf1UfjcBP/n9w7Z6WeWAhSzEmq0KjFV7P8JLtzzzcUqGi9468etifoZBKLu
LkBWd3nfQhj84vbxUoBKf8Y1750aRUVnQ1QApdmIUClCA1TtNfrabNQNCFsAdjTz
wC8cSMA432xJW4Mo5dxzwVJHjh1pNyXJPmp7k5A7pTPNyoK0h2IXvjPEAAeMQglS
xmFnf4iCThj19NmM/DMlP+1XyWNBDCs86+e8lA5oRH8AsHjhJ3qc9yHTcor4sFEQ
+5HftWs57ZY/rhBQy8MKhsJC0Yxw7pOcLMYpAiVoYhQMF4MF7fwyUIG8RAQdUht8
8DPeRygzDSnYeC4ERXatH3sqv4o/PdmvKW5HjgAdrt/Pzf1nmWN236LXD7slbNKm
R8gpExnB+FLPQ6TcaBchG04xURRSar2Z+/aWXNMESUsYlPwV2rvT4R5Ct4NfJycl
1BSuF/BpaDsUB7gOQ9IMYc9pM8vU4B+MzjroIjm5uFLoAHHvAhTh6qCd8UViYMxL
A0L4TsBSmZ2XZfFXm9Oin3ZoZhjq6WEjITb6MUtDX7j34cFnlHygBGjsba8v7e34
IIvVeqE8r8ojUUAE9TVhWh+xNAeHWLfnjNatG7XLm0JkBX1uJy20yL9wpPPkd0Fp
FfxxA3Xh9ns3TQefheqXB+GjFz7IBFhC4dJa8li7Z021Dq3WyBtbiOvzigt6uCcj
wanRGjPjgx8pYTuWbnB2toFBn0TFaDPl5uCW/2R1GqSqQB9ExsPJM267AE3MP3zO
RXPzcZUEgwnnHzpXPD1bd+KQSNY4Ak5wYpdW2d+lFnGI+AgQjEYyWXdpjbVWhmT1
AmSKMAQIcLn/IJemOkxtNEDwvW+lLo2xYfzHbtD5X9jn4Wu1J4Bk8zRM98go648a
EwLA0ZOJw0ZksdDHazFeu3pn0lCB3qjZbjSjCcXEsYJGEmwkx/wWso65PMb5KLCM
F4lhxWS6atqqcicm6a9C9i8TMpR97eqtJTbxfn5KkCCyLFE6w1Nspxv9sllPQEHV
0uZrAj9CCsyM2axmMZ3x13LpE2E045A2awCGN6XD2VpDIt++LckfASQmlCBzk2gg
6aSerkBIiy9ythJcTt5Ydd2XMKjtHBDalI1QQUwowQdsPZ5bxPRAB+ORaH2eU0f0
sj+YLViumyHtGaqQUYY3EdRf+Fl2S59Y60HfWkip7L8nImVqOR64CgcDcOKk7k4I
tOo5iGqChw9xtEYkNaYAOq8zl+OIAaePoAuIm3UanKKFzXZAJiBCsTue+qErewN8
y1dKvmjJMCbC66tcqlPogqzASS+wTN9X02yfB61huGroBSTYkjJcLVdF5Cy3kyCm
GPeVY/8Mp+F/AKYmKkwIQXJYAB8Jq2RXEn24Ju8TlJSBK7Yc86PFl4lAmBs+dXSS
nHClhziHvHQBYdvtz8JIZl2jWYdesS50pr+0drpiji9qabJp6EJ3c7Y6OUE+B3rt
dsq+TEFOlk38RSWrCQ+muy0EEnhSroLg6i3LHdO6QCX/o4Xds2TbqxVpXyGny6sg
kdicUsvOWOTrtEqNQRMYQWkkGd6oweUU4fZec9Qnwyefiir71oWpVW8wz5FdT/hU
NstWX2W+ZPwfQSO/gB7gzk1wp0cjxTH+Fhv5dLBJIu9NkKr6ywYBF/6pqiioPh/u
JOVDC55GJvQfzTcDu2o4hW8rCjb6WG1Bkkl7YLt5pqqa934/jMi2ZtMzBhFn+c5n
UxaInNCInlEofv+hhEt4vaRQu5TNYAqqVmwr9BRAmxDHT80Vh8lBE0mG1+r4soVc
42xKURfzUmqCW8GRboFcSjXFCS35Z03fcyYHtktgqAOv46norvkqKmJXIKjTOzWw
uKXKUFwCCQaVdyiyP4Gs2xdDvir1hlnEVcyCrw45/1u802PTb1GR9z98Qnpk4BDv
Boj0BNa6Q9lZqXp+pIdYShlsvZgocMq8epSaQxhnIsHDVcRcu27sMVfYF5H20iqa
vLO0umZ3v/8BXuEUNuX3ggxAaxiNP4swzN4v6RIrBSNqJWvOxMI0Gx+FxcC3/RSu
r402x5/mzG6pXVldkcwvp4BkOWOK2OQyT9SrLttjDqJvw00u0R0AEwxm2muCAKRv
o5OTdBgTFgrF2E74dGyWaBeGNobivaBIGz1V7iLbHX9A5hYwBWGEoxwe/h52fuvs
ZHDPoLh6nlKiM9MTcY7sSqRZqq6cXbbARrf4x0xm19PW23xK0GRQMnzvcNKVLCgZ
lKZumZO4TxVapt9tkac37O2bx0VcutGi5tjvxkPzDFBVJ/wRe74DZ6aSuB/PoGQW
Fh6HSLWEWpZtP2fF/DwTy8QP9PqUAWIL7gZ8xnYOUFGk0WknNURGbQVUEb8f7wXQ
1JmMtfxJ3gKWkODHWgEWjAJX0Phx7+7VA7t9MUvfbqHMsugsDBByJMZg1lvHM3u0
mR9wE92eIaPPRGvssT9pyg2Ou4KIwuGnoCZwpYzXRIDyEDZ7L4DH56UsMwYVwchv
UufGLYVEFeijeK31dfNXtJ+7E0MapkaPZJUvobgyqW2b2zShTZtLOzDSZsmSyFI2
F4yhdOazb7qSXIugf1F0SGaPE7zi6hp9yUC80T9ewbJfDMZWBI90sDLx5o4OgRjm
kglIlK9r7tQyHiF6WLXm3PJMrqY7crY78j1T76rHpOqKlMibJo58aNLmc7WvmsXd
lhNpdJCwBS2HtrNiHBLozqg5Cn3uVGvfyvTCMGOeOj1fF9RUVRS0Q115hAN8kNSm
Xk7TslO2B5qFW0C/OK3HpR0VVj4vDSeEGhS2ozMs/llX+L/LOBx+847gaLenDxNf
x8YrWAxNtnme8vMGjsBTxErehx2QVlwVMQWD5oSP8unswoX3eHKQDzegHnbRkvO8
Hl6iw243qZgbgSI48tNB6uu0G7e2vcRyAAsLxd2vcJOwbZ7wn8mo6IChXqhQ2MNu
BiGMx3ggyEsH9Mg5hc0vWhbpW2Od01LzcdQMGhVLsp0cJ1W+rnICToWRGV4mDd0z
5uL9OFgMv06NWNsw5rSABwGr8P9Fha6wTaQUoS1drM4OTTXQPhhTEaDVmZ03haVN
9jIQ7s6H9gNGNvgqwYsfHOrOTiGOGgPnKHLvMwWMWOpJXwkN7Shqfh4sqDy6NIZT
7GKoODohCHuBKNKTtuwftwOmeAuVxYVR7WBLQs6ZISVQOvJWIvfm2Y+JSOzGz22n
M8tKyh58bQ5G6i0f5xW9CIcGXDXg/cTR4Yl9rCpNU5BLGYSvJ2UBMb9pgIezeG27
H9QgLPcbHPNKxGTzF0/6oYCs3vXCLzZRXdXiGDRgjRqmqyM/fz9RYkQKedUEyRGK
GoXkzAlt/m5QAHId2+hr6OgfpqO6foFg4HYVgSJy8QnRV385rsfy+8sXRdpDLprR
PbA6w9kBXD8ZntgmjqmQpwn9/3j3PZQeMUdJt8BTNctriAeKRSHZucfCnRoxKLgz
VV28XdMS6PceJntjkuoKIlM1dErsGvR5ig2int60eC4VpMDEpWU5X/P/GKKa5CZ0
hG1kJrfMjGa9frm22u5nK/YxeqGbjqE6L32bTNc68B1yYsA6Iq5BlEp/T1e1fDSs
XwIf9XgDW+cCsrDk5QBPpwbd0Y5ycpkIcdFYckL/31FbywfTxZrjXdXYg8trbtri
1qWJj+XpRB6vBkm3IOtVhSdkXQX742bjDTlNgyX1OoeXMbBmgjgnS0sebC9sA7Kn
qGhJ/r1YVfEoUvisdyGY3oIJjXBtTwSqLOkurLBUxxg4mYfPF3T3yCat2v68DnUP
UAEX2vpii0So1SEuiUAdJsrGMJWN4IDjuli1ThKEbnD7mvcdnG/Xqx7EFNhoYKy5
9/y/Uzub0iEbOpi8k9bfjAxxs6xkuKKFisKqtFMQ0Q1zrfBB287W/5/dZ1/1O+4g
kD9hg8K/yx4U1bB5bvJQ/7njS2gMHVQwhaf87JBYUm/yy1Hf2LobEdEHYa7U60Zm
bLwlKhr6swqGNe+pXmWrj7S4HFTpNL8qELq9U2dW2530SjXnmmqkaXTwmu+wfVAG
yts2ihWmy5ckrqLBfWqKNK4jYGkOL9ULnEhPbcqlEpsUPYRh5++ngiMLBGlLz2Gb
4kTu9u+JuRNMlLGyIfHDe+v0RNSb/Xbv/4b7wolvD+ODUCtMcV0M++J3fewyPObT
FB+sc2yehbFYxP8CgFngiVrWev9UojIwEULvwYq0f/YKKdD7IZv63+YFH2m8qiQz
/IfY15Z1j7JADWq1MjWTCJyfZO0P0jzxbA7yWaadSH6V6V3FJW2P7hRFAMj+b8S3
QP/5NN1K936gUNBuoH5Iqj/tfcTY4ub67u/ccqKwFyLGKBqIRRRCW8yy8A5moq7u
MTLjum5YdaVU0x8vAlrCo0dH7GWO/guoQnfqShI6D05VCUXno65feiF0uAprqYkg
tYbh7WeAO8HuApF19aCdcfSe7x0ouZY7AJcKbIFdsg4V+w67OgKYFKm/BUP+70eG
m0oAc+PixBsrYjjOGnM+mq7LGOWeTLLhd+00H6dvcMfhNqIo04psApBHz0A+VjYo
ArA482JvZxmXQ6O25569A9saNp6qLIXrFeQYEEBTRjWMrBXmJhELJLWfqmAKQ1Jg
JKn7l3RL4xeHRXUGNIq2auDYjOjFZukkG7qp9lenP5yW4mAkh9+kGrjw962n2mJF
sfNHDA01GyL7xWtVXUhONorlwwMnqftOWR3xZCDnCiE+voWt9JPTM1a++MfX7pKM
pJbIQWMpZl5Jnl+KXpM94civPYiLqzOxzCWovy+p0XEXgmIGFpESPHyy22gGkpwN
GgTdna5V9XSBDW98fKFknIqq8ObGsbYiiu3ahvUX8T+aceE8xAFSa+cCXvbsparP
ctAXZz38Mexwi/NuD8KmP8NK5PJuYvcojcMgI9E5YV1Pp42hMNwlTJnSNyix9GwO
yUqmkn57SjvG8QapOcFA2b5AtYrC6Kx/9igeuuDqFuryH23iB3H+fXghwynILf5Q
TZ2sDHDWmsFWv8bQtmz7cRIzuPcJXjIJdZSGzUScHnoYBZT7BcoR+PnWz61GG5ON
u9XHmasGXNtG39ffd2befVNau4qrSr1sKkMG8qOgJX/I9+ylhhl6lq4ATgN08n4U
sL5NwiPh3Cq+nycY1QaGKDB9deSCqJcKo7fB0cJvUI81jhYbEEwjDb+nV+g8KnTl
yq9bxgfQZqKPP5aXGRSG9f2774+R+qooWGC4yuEtw3maJPh8UAmJgHMW7rWfCTil
4Wz5DmTcUjUnOQeB5zlZDG6KiDt5Juxc6sk/WRvxxthc/MIxVDXe+p2FF47eKxcM
mHGIzGgHaGq7FHm4+mm+hdAnOym4affMoLoIYvQXpu9X4+TbIqLACwdHSgdg9Kni
xAdt921u2xjbSGXXdgmL1v6+kOgCQT6AcGaWh0YTUk7xJ7uC6v6GidrrCOS7tQ9F
MlNOqFQeWy+FRf5rN+tkAMctDvlXzICyaNUD+WR24C4Ez76jOSht5U9BK0US1Fg0
PXx9Y8/F4lp0jkQxYDpozExdk5gWtDblTjFu1vBcx4YvU9D49f2sHjF+owClw240
8xS8gPNT3z1d/ahl1wtzRrYM1iHr4bivr6wsE7Np4rajShhVnz8hpYyV5Nbzl0UG
R/YZQESkcCuc+jXualmLZ9gqzvdmT70pfc4fiTOIfJklXxNiDoxZbeKrOV4qjASO
T+F+1BFlPPtUgSLBtSTt41F6orfn6GgNiOGBThVpuQ3lqjK/Bq/5Z9mjeGv48nMZ
ScYOrbedC+SUAAY9Sb3lAB5OQUHOgrG799lVEqQmzLWQHGYuIa9RnNgh5Z7nC6YC
BpfZl9up5vstdRL8dXkEk34K/4dBP2tzQ+i+0w/TME9mxXdev0rUUAaB4A+pi9UX
d7I8kEa9MT1j/0a4RQETgVF5g5wd7lhBiuL1zJKTa/A77M0b5zBHugF5tfPSUExY
GL6APG5B219YCnpaTmxVtxc4hIUMxytw7Rd7EvKfKJgJ3ovKhEqmrLdlQN3sLJRZ
NB4x/hPBtyUUduo80sb2O7uQAhtQZlGc/0OR9oFnVVi19GY2DT7zy7XeWLf+TDot
jhsGDdTmvRypWfPXF6ld/DNasAHGlqlu9qQ1vCxvqHyzuoytF3TYYQ1swzSURzDn
LdsZUl3zJ2aeahomLf3bsg7+ux8m3sOJt/o2jgTN4JBrQkzP0Z5Vxi+9R0lt/QVV
QyXlNGHSrqo2YmtqdpS9gQOnNn69vm4U2tEf20mc/8JzroOMpgjXjJGNyAGqgVYD
SUiPD8UmV7Ji1pXkCKWWymgwSrWPhmmu5wSyOWeZQQ37X30zFplvmaRQMiWVqlIT
Vw56MqsrIOv6z2FeqxlgsW93QLVlYJA8+UQI1DUQk1VFhofKNJL8kqSqLkLg9VGe
03EK47FsoSDdo34clu9KbwggnKn/jyfi/bYTjfjckWzRZPAe0lfmNkbXHN1xGQQM
JJSO9lHE7H4Le0RNSfXw9UV8qeqpcyI11YBj5kypJhef65vIsZECNS3H4EE07yqM
BuELn8ZW42F7jfxcecg8PPXkxN0tiMJeUW412gV7Mj+Sw3armrmkYFiB03ZRHJY9
SfC1dZQ+s+HC1ImMUMfrGu4x65YAGnGuBjJ5AdWSo+iGSEPXim/56FzCm2BVxWBQ
XJyyFmmGhKx+IffgwPkt0bpK3XjgywN0JfuiS3vSKKgLJC2zsewcgUDm50kgFXjX
1IHA9L9/4R19hwNGKK0CQ3F4/BzWZzd9RlJYeiq2VMLc+4J1yw7oTQVEk1pj1hBB
3Kos5qctVlpf4YEQFjwkoX2HShAj9C45AgQEeCaecmH6js2hZRkHF70wo4K/HdIY
+M0V2oSX+WL5AFfk/ViLxqgbhwOetcMoPoOJ26tdTMFyDgBjmTQicjoFYoSLNLRE
I0lTHH/W91F4XeWPoGNLiS3vybSZiDqTKSBZeUHoNJmhcn9CWKOtl4ilvrZNalqU
9B7TQnS4GVJtC1vQak8AU9O87mT5hBcNqSAAu1yiop0yl+r3c0vxZg5Dd0OgN2yC
ln/NhByxDAN5iBTa4tnBTX18Hq3gUyHobv50bJ6gGuPXnHJW7K6SehuRZnKa0krt
g60wC2f4sd9G2RA2RSC1uyHOqoVnxOHEEuOAF6vldhdpX27B6X+OVtlpizdEu++Q
WMjRN6ua18mCGBP/YEWorEYoY/thg7mldW4HqXrzEecUogc+5CjOm1HYFYGikdF+
50UIaZ874lARYub891255K16EspdcXRmaARjWCSD1pZqr6vE7HyT1fXViSuUln6N
EFOlD0sYBgsmlOUuh70KXcB9rGTIeH8Yw0ukek4lPg6AIvbsSAl0fRbeGghVot4F
3NG+v6dx6Bmci0xsEECEXISdm0Nim4c/vZlNyLuEOGGqgvgvl5dVqb31cXmykUS2
TYHH7DeMaKkk0/26Nt92GUen6+nPiSZl2o8yqzy3SEQw/TW6S5DGELkCgTotYsFX
3zKJJS78+hMY6V3mwDZJABhaA7wfi0rUJgmobEIU0aN0elE75HtQ9MFt9GKPtU68
6TpF2uLIHyNoFL9ulqps2AW25jkfU0+ObkoFUhsiBrhdAi1jAtZzmIMrpshcgylL
0fgC/VkBGseuGSWS6KCMyVUJGicYzukfGa9lhxxIrY1GvKYQJVNC+HUcb+sAvCYB
7nfbGBlAnUHwW9HOu6+j5E2zNfVUvnwEEBeP3Lee8TMYunVBM7Xx7Okyo+75C8B6
T+///JaduixW4AMdo2LbHcJL2dym6Z98eeeO9K/lsLvToNGGbKs1/8SXzqbONiWQ
xb3PCgte4aa6e7Onas+axAUb/T3VbY8x3oYTlcS4SPhIoC/xIe8b07b9i/+0RHWR
NcXeCA/hd5VtHEd+f6O53jfIzm5X+rUyDEWvAe2ixQ5neJ10LQmeZJGinBgX7bxB
+I8rF6VQc6VCIRTGo6noqxGS74YLsbsKXONvU60IfbTGHn3oAlikySXCsJQORGGl
T66GCGnO0uQHjUympduiwpNbc8KS6JDHSLq9AphPxnucH60VEbPYDlOOFBYBdJvL
d2Y7MJwsdyOwpt55FocZlbvEO0CxE0VUIce1+8rT6pwTq5/m3xg574VDXSXdlPj2
Vu9Iv7Xh4RudQyUhrqmqOOftGw8JCFANRHjGxIMB+lBt9j8G6ZSeW3X1hdjRJig2
FQybQqmBxcpiCpHN+/y8rrtH2fUCXcyHk6ll0BQqEM1SiqYTiw+/IxsPxkmDhkKS
s1GhQrTvxBRkK8v0BkSQC15X1gG9zXlfDbqyeH04WxaUizGStfwfQiy62OjAFnh2
8iPi4SIniHE6DQLMSsW4wOgPWhRDNnH05Pcb17nch+Pr47W7n+fWQYf8qxoCfy9y
l6dKm2R0Yv+kjJIYBPN3nBe0l74/zOl1pliFklHDXN5j1KeNOGAyCPIWB9AUmrza
tMejR10cxQtl9cl4nt2uiZls75y3+vxO8YJ4ApFX1ss1CDWeDTd+fNKrHKy+ul/H
4B02IKVtERKQaw3YMna7rCIAO/DXyEssbBCYiP3u7ZIy4Q7Frpb6BV2BLvodKps3
vFk/hW38Bc+y7bO+goy3kJIklnxPtobNdGtw465I/YZub1gAd2qFrO2hkg+8cJug
OOo2J4KQqW2StaQ7Bj4YKxm9/cg6RcyqjX/pUFdRThUrubx17I6NzFHFVzUKIN/b
Q9FFWlqiBOrYmvfNEmzSGITKZrsuyNuHmG3ZR/WNBCpFd6+IKBMKzhk9Ijoz598B
qA1aqzhbXHPHkxeX9HgI6dyUgrXj1PAxisSVUDfuwzczX2WcbgtWWYUFaOKlKhaa
35KEQEvUHGem9JuY5B/ZdQ2D4vBbmpukRLpEng6YDNxH3fy2WMz6JaiDZLNaow/W
QllAJcWrczTgb1oMGKuTEvg8XQybeXS6ziUCTp/wweWB8eAQV/Trzk2/41z1yWUh
GExN72hR4FSXWtGHRzfIVajZeGRXJPqlhD9zkEgn9PsJQ1GLq7WkzA70nJo2vvoK
QKcS/Loev3nPDmfgf7H+5v5TXYzmnoNmmTtoa1zCWmLaKEt3v6GtvjAgv1mz1LCZ
addDvMz3vI0AtT0GIoyFdogpWGYVWW2UKVObs7UUXdjTXqoQpzzwTo84COjwp7hR
hclMdIY97TcsSRg5Lz0lRHCXuO4OKobJYBGXyygUv3fbtY/PeIxVm8QSkKXeRWlI
WnkP734A6Ad1h9tCsIy+WiYpam+2lVuO39lx1rwv4bwQTUikSrrWPyvIC5eOsHh1
zW/58qpCfX/ULPlx2pW7ZkR3clGQojvhxBjm/nfnKbPHc2epy9juaAI11/R+UITR
teTHBVSIQ7/sN1A03I6c7SlkckrpDZ/HZPqNL8Wm9qS91sytz9GJaBz7wufcxIXv
8GHOaQgON2UXDzKFG5TdqBhzC8ttKIAnkgiK9x2Ir7BGlQCM8Mv/azyccfUOK1nX
x2i7J0jXTc09Rk8DHaxMdz8qi5XEnXzrsOQa5EvMaXtPeXHNxH+9JKzi3aXy5mW8
s//dpTeH96k+FdQWP1pORNxMe0Rlqdt74vSkceH3h6oCo913LjISXQGGFoEtAVmC
zVq5o5DxvWko9p+LFdL1ZO7jODLsWvX/VWBEDmj0wA4G/zjj3sLzdGCtB6HEqU1C
3WXr4oDXw/v+ICOtNsKNmNMvJTmwSbBT8YvjudCHTxQzWEwBCeFJdE+d6eYVTLBT
Rs6gHabdPjVRAjWzKlaXkV8eUUH0YWNGOhUycwh/ppjwZnfm4M9PcgUMrKkVJPUa
uwiC8RTkO/BQuLaI3syGgGGgsw7N289BWm4/Ocoe6AbT4CLn9cFZjg9w2AOZKxtN
G4doHwirHZKLQyIKMHYZ/TILKsdFxFOI/fANq9G++eZRq4aLHmOXKCUCecWXH3Dk
G11PAqDvkuggh5V3qbl739vVevWGjf3ww79MSbAUU8ja/YBCUPljyr/vIoB8f6Oy
aemYsyElU0vjI+fFixqpd0qJnzuHOhpH/vlFTSl8n5J0CECdS19nXhUaaP+o8des
ILoKntRazH0Sn3FrGJ2B90YBzfAXghkqdcp//CFUO7YV46bMSzp3QLsz4lmXdx6z
lojn0Xa9dYvp2G5Cq/4gOL9MLWtdxXPzgWogaAXe60AP9o91hsJjXvt6P8jVM4BC
bL8dds+N1lpI5lqCrrl8CT9B7yZqQ8aiBz0OxOe9jOaa+n0V3IznQhSmg15PTzfO
NuCiXyoE2q0zkuIcUFU2YouRa8FIWa5UoF9Zp/rlJuC4dcz2cObcuuBVz7wZ3CCN
lREN+PbZX/jP58vvbB7drfjfof8hJtSYHxet4UUvT0Jy12d/kHvLCDUTOQ5dvWya
b1ge6w9NyohfKfO6i49172qYN3Px0ha9ujQVvGDXA5YTQ1ATV/b/5MGddb1Ia/gq
aJl/BbQrmoF6sQiK+ZheHYLSZWd1wff2681U+UN15aNacveCsTgWtgR+6vHNaEWy
hRqrbEyFzoZYSCf407vkCvEJMwjnmQdCNfWx6bQqqEgYRH/GX/pTMo2TpSpG21mF
6+qtL1SleQQ0XVVSJauhDTx5rmzrIsfXfAjfKR1K01cITv67tJh70+iajnO8JUOD
uGC3C4yA29H43A5KpTNkp0/bR8cRwDv3EqCpLCOTXQA5fVhpSOG5Z8Ub2k0ZBeww
5oumLvmO2polQ+8cJqJZqMyl9maFc1Im3plIIWKjBHE+RTYgOvw5yj01yNjWDafB
t6ITQXAW28E9uUAvr6N7L3Xjn/jdbOktgUB085AQkab31jZmLQ2ZbycQmaER7rjJ
IBgBCewQfBwzLxdb7xaLnY3OKMIKye6FVA0yqt0qMJ/42aHxcYqOgrNKDi/LqlDH
/E3MSSGdWM+WGA+LPX21W1NCJITT+ehAorefQVYP447vUV/GbBMdt+GZjGKYMWx0
7yVeHSbXfxGoFndqHFdH9hLC8PxmgHMZfxfDdyyRGvzKAeo4H3JWyfTBkHDuSptN
ln99Epg+HueSSQr+m0R6z5UavBM1m//JLGS34+9B23cLN438akgQt6yT7dlXQ1bK
eKzGSWQZqBExatKi8qSU5sR3B5vMpe2wD2UHWPDCVGtGrIAOEZvVYTcAN1hRavvW
9nOvWZFQsr9U98jUXPQL/591aizUCDSRTPoRCl8Yr8WoyK0gh5YMdmbuXE0MU3D0
c5j2V/aL64GwPB8FgL/lFgClKEDx0Z3AvA2fMsa5bidqReqkmzz96qZejrlV0H/C
GUll9yYyavzPezRvjxvx9OUfEzJe634dMiwbGxSsQv0b03YI6KecMC0Jgw6gMW4P
NCsW5/3hpH6jpgrCFSeiir376BL2TgjVpGXxx+5v4I/JwUgQQ/+vMA2LQbU4YbbU
fFCjsodoLvaVfjbQnORkqW3Elw0IEP4gUVG1gpVt0XMFxv9u9dlhubc8TUWJNOLO
7aJbtFLXHcr/2H+nnexMKhA5ImkqxuoUnGFpFvd8BEeDpSV6a2bvwua20lWSa6Is
+g/ewGiZOefpo8zo6ToIn2wm4fMegPQ462cWhH0WWnE3bmVzECH7jMuChWrB78Ic
SR1T4sNFiLWj88x1kotelJABsq4/c1Njjs3g8cn5rJ9M28VdA4XZFablxjTXvVU4
WmQUj+xUfSCiBM2zGssX653gDuzEsWcqbDuTmU2fmX0YDhoiWWDCK/vaI9Ynk8aJ
lE/PUrO8MNmyghmQVkVJokfTmN3RqC0RD5+WvHljlajquK/2b3jDXAl3oIag3mpr
2ABt/2FLAtUFqymtoNUqMhSY8Pd1gM4rrkOqnK+NjKaW/EOdmxa3i/f4OPgP1Jr5
i4oj4KpdUc1fDAkBVqigb+dABxnYMz1+dt6M1aawHGPzit9EtXwC9cP/kEnaSBy0
n7I2XV+Z7YKZQsEtJAgBfV3zEqd4INEzPBblSQLiePZYINll+oMHzIeMRts28p7h
/lknmX3tZ59Hepeu4DQLRQMH+RIVAV0xx89Dbk6kiZFb6BAON9Y33gfd1lbJDpZU
yVxJyQ5F9d6QRUT+on5BiIkyydL6UIp7Ntv8qEAz/mEiAg9gsUkAPue/Uem5n4s5
OaISeJYxmMBTSrpTjyrVxz3amNZ8+jp8D20rep5MXlfAB+f8aEUtT8fCvM0W4Fsw
Au30gL12u7g3HHwBCgi2N+zz3JjOJce1vfNyfmE+1F6fIRqpoem2YHGlvmt1/JGf
3YM4geAqjzjv5vwnYaiQErkRNIY1oHquc1ppnJts2lQNgscLh0S/p+Bt1dy9YNLR
cxFVGXfFeiGQca6PhDmV8uzes7/bq7Cv3lspZNYMiFjnRyOw5e2medQjiToBVhEl
ExRnD7lSeqk8D42XUmXgnsEGNS5koZ0KgcK+Pwu8FbUabg+Z1fTmt/TqjdRh5Gpo
gcDIuVME4NfdXqIIADt5EZbqi8XpHvIePJkYXj5KigAsXwXjgbrG+/G8EsBo29Tr
xNLO3jhRSMRGfIDLqkRF2TTYtuspT4/sZEa3yf1AOHWHwNkoDBuWWsnsP4u0pl5L
F5uwD4ORZosYB4msCNPfIb9Iu2lNQMt6O/uewiXXfFafXf0YNjC5YTMqEkrnLK80
HlcVvnJXZh71RTsANjSSsdBS5wI8BNFgHOG/4+BOuxN3OzulFAvQfqLYmKvULDqJ
c9bIC7lVDg3g/N7uWAykrT9/rZcGpVXomMcMEd186E4b04MXEAw1Q2ZjIaw+F1cr
+HCbCycOQgna+jEWu4+yXUBZV8ZXIWdsq7GStLCLjNd/dKHIWJsXaiOUY2G9xPOx
AzQ7gc2blRnibzDmVDqzQEqcPsoBEHKUl1TD0YyGJ6HsfnRk8vh2Sg0Yq/tjmOEr
qa9AhI+YJxHmFcM8KuZXwgONeAJ/0hMMPn/YX2tAFcO92PT2tyECQEQkFquUH/8K
aCtpQpXq76XOLpCNL8fOI2f3pcQsmzhu7Pl+Cd1hePfbXDGK2TjItuBsU+xgyF6W
nw5dQ4GuhIWk1sAE1CFgh8sz6vHAmRmLZvne9UDR+In1oCJSq2RfGlUI2N1SXn1I
iHZ2gefob8VNa3KY3KuHMXEXy7zPcrjgH5z02AgAzJl0SSR/ni9hE1BeA378wq/q
C2oO1GXqYTV6g/btJWUWwbE8sAixZDtO1JUvDBsVIjmqkJW3+UHohTehCRrF70ra
7pwrJExFZCqfwfAwl6CWEwCUnDTb9q1pkXp7NvUMt21UqHt1g5uiNqq4GXdRpRCH
9OSO4n/5smvdZnvIYJFq1VKKDL7IdupUqr24J4RUUe/FlwsuSVpJDruGbDZ94VDd
NGkxAZdQjR+s+SvPzTOX2gt0ilgOCzM9UzZISDKy/1HikpnJBwYr+0KhfeIrAFMN
io/S94KwW7FfusrBAWB7T2v0IGnIxNz5lT8Po/1EAJ1HU5lN4Z41IYaPTbL2Fcnn
KGcJvlb5/PS6wLxGBqB7zK/MZbU4TXcTsAddeDS8611VA6m7RwctpyeTkz7W2Na1
zwnia9ciWcWt19EZAqFHqzgoXfB36Yb52y9AXOlTouemvqBnJ8UWLRek1dYmk8F2
ghPLnaMAYS45P591DTOAP4znUx5cgFsfPbnqVzL0QjFC3Y96fQVc/DZRpuha3i9b
G/7kgU17yAqiIPj4nD6H5vMh5w3i7S1jV90UfUbjhqwas5YiLa3unBJQA2JUN54/
H8loAiuGP4aJrsi2Ffa2N8LjTAGF1/IxO9b6FxLDfNmWgzVNC1wQiCu99uXz8XzA
hA8PYm6njwimpTmJLkx15v1T2BvWT6z3ZXMudk6m8aCCAgJ5I/vLBeA3hDWU8AJi
Fu4sooqSiKvoxK+2B2AKoHMaJGD6ZkrP8WkFqHc2EhsFMs4N54L8apzlXFYPjmdt
GhJS3Y1CtPZz8OJtehLdkXbAUkCfAgBdjooh3N1EcJ865QKWaM/qkodbTs9vPlq4
tGQzVqanmtrkGTajTzavWvLTd1b71jwIjnOGFLU3FvHnjKwdol0+u4MaI3Yvuskn
PFelZEiZSA1bUlKynUPzoq3Zr/MkoRdmGYB1eHmi1PYKD1yV3xIpqt4eyscYnLW9
ZtLAkoLsKGTg3u8RQXDZKUzSs7uMJF65gPSP1IkFZWIx1SxUdngjTkgKqjG11Vkx
apBi1d/Dm5P7evLd65QF75mhkjSbX2bt9W/oe7iWJnQCq6FFkhCh1fF4uGJdb0R5
XNpnP1ivpMCqbUsvFRFFGCosh1Qp3OejPKM4cAjO7MUEe2gUvYjHM2/s7FJGXYXX
R/st4kS6tp+/rTrOrPSPN3SQwuRMyPdULG9KjxwfLjM/U7m4WWVFcAWLTcSoamGg
BcwaphDqFnclaeKJyx/p1l651RHLl1qHHjf7Tj6GpU6vAw/dVwlGi//Bk7sQCVcI
gLM31ukv5Ogs8XS+d4dTySAx4zqkf8FlaHg9VZd/76QTbGtAbzP8H/ucrftH3Us4
0krFl/GMgIC1athOniNgv0xp8qfL73fdu0LZGnDrkgZLjhZMTcNOpCk62rDQl7BE
TFf6yvszRQAoFiOxXPRjIrQD7JG2salSXtht7dtL6Wf33CGqWq3LZFg5dSBe3IBU
kybcqDAn5Z4O2Yt55LV0G7/RwfNDwjdtmhmpcC5q+g2UfOrzenfl0Z1zeT00cjC4
VpfPMkkar+bJMx/H+mO2fwDbG6LOwAh37AFrqRReFGHbxcw0eId1by7xU1rRWjGA
x5QdO1RE4Frr/vEcP7nMx/m8/hxBE5u1Ysr0KFrKK/lt5oLcbLBC2/dO6P8VQRa9
x/cxMDZ46ISq5iCCX/v7IPsaBglafc9jSKxQ0r6PL0qs84GcPHNZURQwSeggn3sO
6zFDqbrkogxLG20V6DI98XbXatyckaa2BQ60LLpIxtNIl+171JyHQfDwQHEMWkej
RVLXNtVBe4Tf6LZYJJ/nIdgVWuYn0wprXOT97MPUOhJ66MD2TXLGgt8xZ/rAhvQx
PAVmof34UmMlwGfHuZBNZSgQP7M1wW/h2GZ0XLqZqWGp/zQPMLGwUS07SnAgf8S2
q3me0smq3Sk5nqq4r7slUBiovgFXIU5zsED+VZ1tdvFxadVIdNLenM4N/yG7mAMP
jxNx3R7EgsRzhmUgDgTwwlZg6Kiz3PUyYXGKAcbWARH+rto3It3mowEwv+i903X8
c+y1nTiK4cJoiWX6Si19p9Mc9BOUG/kWIl2vh1NmKRS5PXVoTlxRF2klq8sI05I5
tBZvoXZflVHwPxQnd8bMkEgyYFBEab3zwqvMEgfLwgn6njoYRro604bbOKe/eNH0
rYpuHj0cqc+O5dzQtfRwx0z3KXU6ayTvzpidRPqhkaEauySXCPVT1g2XfYlQyDUy
r+Gukr4RIgwBh2dCpc7aVNp2FnsD4fjYmbckDG5x0bpLeoIHXoryUqhOUDQbbKAq
wffdAwXU3nJbH14r4pMf5YFtpUyYozyWgN+cPqcMEauO6P3F4OVRvGuFYsEEo4W5
aX1qX4ubyflClxJJjL6b2sPwnK7L89BEpmHLMQOfyYsciuKJVP8rAEdevIFUUtsL
Nd+tZQz2c0hlGXdWkObTDMpAjBfS2UXuhYVXJiBxaSpi4fZNnMmJ685evBTg5A7U
kZaMurNVUNKaJhdAMhIXoxyn0ZHTDxYQB40vGxdKgO1fnVs0h8SIrkenKm60wREY
ByIvmihTGyC8/R33F/koL3qcI45xuB/qEz73lnOLfaPmtQ5rMOJVmZCvxsxdLrVA
TO/kZPVPBk9K55nJGnIVvG78dG4xQz/o5M2Cs3MTlmdixFaMT1JUQpJNpNPqnWLL
sR3QD003hEKhHPR6bKJf7aIlGz0wToTaJ0+VFpvmNAxRuQd6LWb2n6nlNedwb0yY
cyz4J4D7c9lm3U/dt7GMu02a7Nn775OAVxdvDiYoOARx3xf1gjenRtN1j1/INiKz
F76S33FPXjwMe107CoHeZmtpbKsj9oBQvdyox/NHAdow8Js1fiME6RMVBVtbbaX+
BUeC+aDpbOL2BhTLe+oeZqVhdfO6Xf6FQ3ozXquPPqtOrmOdvbD0urnuY0qoTPeX
iyiyBWfFedfwYnaHaMB4h9TQEevdfQkrh0ktk5OQXQv1EkvZCHU08WY/kpNrRsKm
cvRHqBk57kzIqpX055NRbEq3v3QyGL6nGigssbS9oA4mpXFWyfeOUGYm7634CO/m
RNzffQhUt5lG/vZjCpf6uhjzjUOcx9hTjIpTf3nX2QG/usRWoNXq1jqJx6NcCKUt
eVfjAQJ5YIDrNBBfbYoApu91Jlxs+JH69bhcUjrBZZQq8A1UQfcjkdgc++8rNQxa
b10ApOvchOEpHSPwHvy1l6u9VG63d35NwWMSU3Ii2CkX/ZbtQdLfb973VFJi0isd
mP1VFXNX0BiGUP8ypAmFHMBuqmx5mXcfZu8AtoiDcOBIKZ96h40jGCXD/SgbVNJ9
o2baHX3gGh49TQ+VacZBhvZzcOV7ZqfoOMb9c9KxFg33i+24T2NlIZ5hyO83qvTh
KyVruYkcBLkAOIWbfS3O3H44gilVJirAlw+yNljeZNiqdzEkUW7IGwGtQP7trmDL
+uZw1r7srZV2Ow+KvMMQVDVaoJ+7Uerp53sm+pHSCPZ7PiLmh3Br64Xc1LdQor3m
myJ3cVqfKiEtBMKq7+mN/iobaSNZ+6mAjt9jwbgQ2jb/TerUJYs+LRHqUDhoveXJ
YU2KiDEQCVRHqlUEFllIE/Vp06YrAB+pV5wTB6mt/krP4aPatqLZ3PZH89fWBKuV
LPFyV6JDgF6/lbmAckSelX4UHAun3kSYHervbrHn1S2HdYJC4FsUlj7W3lQdwLlj
BHyliXANv8sfRpdL/eNxJYB7EQiNxPgadXBOFXNwknazo/VBlhIDTzfS8i5lxcy9
NLaIpgLC6yVCdLZzR7osuZZA/Rc5NORtfZDepSL6QqrhZlCzWTdtBpQlh7fh5Nfk
N6//btTECjmILyuja6t+GIFrVfaPWbi7DxlALckwbTlB3IHjOvfTa+ju8V1hDwPC
Ob02rGNnC85nvF1W6+gf2Gq9fmrcUjCvD2quWkMafaIwG1BeNRhVWi4Jhu/FO6kM
ei+Rux3iQ7fikiPpkJ7VbikNUoSuDruSdDgDZKW+IjvqryMtCHHH+DFqrHHnAkWj
g2L5sgbI/AFaqbvzxk2lmQ4rLvbd2xHkGe0ST3AlqtqVvlIsGvVC0zMe8yVfkf0V
yJWaYzaC/bXZvPqfQC1X7ypJZ2nq5Uh+WNd/w+HRpQyoe1PwF1Em+vm/j1X2aQvn
oG9w5zmBOW+sVn+qPDJ6A/ibhGzdFk5fTlnQo8sRMzJtST9vN/AVB2/f0r6zovyo
3m8Pa86JndhKA3tjHnPhP4OlUg+cgqUG7/LKdyPECP8jH0eY0K+hQxx3BhXgOwTv
XTHELSEuIZqaiquA4yWhb5y0qKLTI9if9SXcpwvwLlWrmR66gmCyBas5ghLjAcPg
uqggF+jMBLvT8l3bV0L1gypwgPnWf+iIA31fDjZsFBqMu5cKS3XE9DNwcNx1ZJUO
4hK88NC7OTNS1oEf5yRCKmhYsWvKD3ys9dSGSdhr6KF1A4lEDCztPPRcA6iWnEIr
CMkjXx5FvRGLlaO71hTEqwVGmNpPeWbP40wanH5VqcUK7Mhloa3VslBUO1sjLV7/
WEzmfdgzlxsG4weOJ7WH67+zkrEW2tGjjj1OCV0Hpub/mgOks7FqWQSCvgZ73K+/
mVL3mInGkyOdy3VZ6XG63Uv2oeYY93/sIgF47qAT3loZkP1955yqRx5M8LMzb/7Z
GiakKgJAiGY+xzJioIABO+DWUyb3pi1u68gR9e/HWR1YGb3meWjiX3TPwP9PtwZe
wFfuOOV/qFGBNpdPqgV7yfXGJQZ8GVVByFFdSa3rIpGABL+x2AdcmzARaKt5L1ia
pT/bPqxZR21Ynrm3gkBTWjb+/zlFX0cykS/NxYTPzxewM9/Clv7D4uii0uIG5pf4
okXR9eKYQoAzKksnzO4Ci7ux0/dH8oyB0eXFHy3XXQp9MSprGPV4UJoIUW/tKcSS
DI0ZahNVOHe/cddirjaP9Gz0YdCahkkAf7JdywU8f5uWeU5k/OtPGjz9xfdOxqzs
3VXdrBiQjbxseeWOS0GRMGzPGfo0BeP0WA2mLIadDL4HaXS2O1yw7XGTp7hKXIeB
MRYJZLZtswI94Caw2G94Bz84ghsVTO1c2y78DOnxRVLdmY1Q9d5o5g7W4Tybjdau
aBTQD3kgnWnO0XpPnWNX/Sv1xE8hq2n76DwvYgBHtt5KEl5YoRUODT9CbmxvGxw7
//MtOaquT/A7uPbH9BwmUTVVSJcbp7gn2Fti0YrdshukO6jgcImqjF/7cZ67HEUc
Uq/iImQ7Uoz4bwiJ2VTG4DJ+DV/AmO8VOwFWdH5tzkogIJ5OzvJc8JfA5SDerplU
ahnK/4Q+GzAhT7R3L8sy/ppuxWQl7Cs6AXkDci4bayXGFJX36C0698Swac1LgPCf
ToAA0DLfJ/7O1PLiojRINbMG44F7UboveWNNi7QmViVQ4kmyP/l+G1kDKx7LJIdL
1b/zRgCwL0fNEBosjbETmypVu7sli+H1Hwe29g1prIalmM1jMWlofYrxnxygf+fn
iLUwD0HOMdEbUzK/WjbRYcpmdVj+SwvXnWJ8FDouagPmbdPXzdcTMQeIlo7jrc+k
6DBOlKu7HThqYM/Hu3hkWs0Z+cjt3oB3GaTrAQI//bJoC8D6Q+TajYdCIUu+E57l
GmxxOq/fM7RrYjf5jGvYGgHxoJDENgZ+j31WQvnDoh0FddtD1gsAz0JmT2HTG0Bp
DBvoUewZEaqmbLXs6saaPclKFgdCAyIi6srQEEmiTq3PW/zKJ/dpDOhWWBGHHKFr
gOX9DiZuUyBPQNUxbN1wn01LTO+NgWXA9rXaKTDn4BuIk2nbBvt10UAZoqdCAKsi
ZN2pODnqTlW0NDhNCDyIg3pfTYvy9jWGmgCuwPpg+TYYHWQEEEF9crcI8ijUBr6J
2Atf9bLLdGA1Gqdko056Z20QTm4jymKYVaLFxK0OpouZhp8ErJtprAKYonIMwn2c
FzOS+s2WRYgBhih2r876CI6C3CpeVjLz/Gtg97ycCYjXRySU2QQKWOfpfJzXUFDL
dewuQO8TR3NnbJeKfzLStyjAcZlY9mn78wr6vxbqUBCanvh16OwkPAgBhaV0fwN4
O/Ws8VeTl5E3cR99mj1a5JtpVfsnMcPmYaCk5elm1LIaw3yywz43Deuo2J3esSoO
V8iIh2VS+heFY5cM5WPrWxfx6uNF6xUJx99W9wc48pjSQnPJr7agfU/Eqh8MiRx2
Vj+HB+jqFn7K0Lm91x8ZpANUDco9uhKWVULVMRwENAEFe9AGPQM3g+l/ZeBBdv6p
N+HEnQ9TXtC77YJuZI9BcHiX34F3bPxSRZTWB31ZwvXWOGybVyo2PmX/wIzztF1I
eu39ChRnbzjwEgulrAx5FE/fk/XIUObLVn1yKvHb9USxZiYkeEuP1Jsso6drpPOL
e+YpuHL2URv55mREYSGYxT/8gHP+um/6Ojg+4ue1F+jho9M6lC2s0JimHBqFvHqG
pPKmPIt+LbE+Yr8M+yLfPfv+oh6B4F3BiqW+1ByQU/7H98V1Tzd+QtkirwJFnnKe
w3zpdO07hLMwdTo0gSeXfAkvA8l407GPuYW7x30l1nLN66puYC3F0EDR350dYFvF
aVDCuEY0BxHMSBnTzQiPoQztKKzrdwBTH5ib+RQqL3oQ1kSfaNVOCbPI5g4lIGXr
K0mOS7DDWRtHK/Gvwuh+WsWoJryCCuyNTzd1ldgUQeg2au4xHgeokCjb8i58MKk4
u73R5H1W4u6T5wCmHqYjnDSqiyHfHBvxATHYboaO8tsakGuWpFWvzx+KySTcB3m9
3edTlbiQ2yga9LmewONVgJNJ7DpBvYjZH6BZEKM9oM5b/c2sRPecYr30pI6GKjDC
mnn4QXDpuhxONkyrK9GIGp+z/CmnEQfNuiGE2BBveBK+2bxgn6YDErSKgG8U3IPN
kJ07UVjtFQANM9sNYdLq4dQzzUYFSkHBTYusVS7u6vdgp6LzsImy2he+sLjlnfUh
pxhRX+v55xaQ7dwLNLqFjOqKt93R0vZE6j+Oolahu0FH0zGdYnA1tfJ5CcWb7idz
iN0b+9xs6c7KpsmbdDKu4d+BNbG7yLpTSsGKjGx77MRfOp50ibJiy3ywvIwy/1Dr
7LZWolDAC35vJ+eTIE/t+a+KuHDzO210+FCtcL5iT0KXjpnloUkCzqawPXJK01LB
2ZTJv+X56vnRvYH9Q9zVZk7rVLAgi6EbQuMylq4RcVtR8RNOIQNRXv4b81L8Iexe
34/p11zuZj6qX6zHxHCNz1PfIquvKEUG8S1P1uEZR0cY7ZmZh8BWKU8X/Xq0+nuV
zd9Pn3ElKGAieRn3Q/M7BGuL5YSisuH1nerCqVJijZxLdc+ATGMSTosnARJsNhC0
31Pls78plQ86hfO9Nb7QaOkuzWyv48z/wq+wOwyJGvrF6gFVWmi1R1YOSqLQ9SML
N4aBOD4N20vX6oJn6bKzdK2GaS5hBxrychHzR54sxwIwSROvqwQl3yeM9M5xMGr+
ugGFfm2vqa5aS8LC1aLTVp6jh/Ri4LqisjXGz5hhxt962ZW5IjNilFtJ/bRnRucy
eOngLot4hO7UKSCKnOvGUcnwVPYuhYzRbM7Z3RJbRDxsmt+f3MtSXYMdUe+HZQ43
KjNfGkadwkbxAYb2/7sOHePMIeLJkhc5fgl4MJ2EFqlBckNsAcHQm2eJE/50Lpu0
lgGWI+1QM94BjdMUG1F9POpFCNlRzxOzviZYrfUyOodAq4HW2H6VHm5/s6sU6d24
7yXIXkXsKh5dU4mbXYZk2SvJUwor+5GAnQAmKC5hXteVSaXxwxJ71aafXHEutoOF
npK84DiiIhuUYIRTln1+UwnSpG8R437xdcdWfclsmCKXm5bKvC+z+BfWAqF4MduT
M2t+Q6cDiSP30GqVcIVaIy7cAAlNfXfzuCw1QBS9Hu3Q+pONq67FY2UipYgamwzn
eGQ+dGn+s977UUeYucpYqP40Ct5aM6qI2INtF7kMxdAB4QeaeH9sjGANQqHcJA8L
Hr25Dwb/jtYwF7ISHoOocQqCZ3Q1W/swYCwlzf1Xz4sURNoEyX7/ioVfUoPy/Z4J
zLQqnJKeJbkMuDKlqV6+0WD/MNJp4q48chYQ5LaYHRPPk7sjikVIzIrKKRIpyWji
IfSedNuGSHZahduOOOmAlQm+lQeIBSrHWbxim3whvjZke2mLOTwgco2eEW76eQia
L13O/im9ESiSxLpm0EGHOm8MENLimrrlj9lx8SwzviuqKIpZ69Sb7Q0ux4i5rvEg
Mco9qyfMfVfAnIzcFnUuxsa9dIPc/9j3pJrh6uBdtSgpR7+fEdpXQgncnBCCDVpi
WvlKdTnHWhodBhxss9sH2libBd7D0Jk58xGjvy14vxYK9vDmJEXuhNIP0otv4dkY
/FV/QoB46HQtT2Hw1RJup78ZDsSVLXh7h6I5oBcoUuIMbntASghPbYE7GlhUM1iR
nAS0pT5lxbBK/szrFEw+odojzTCNg0eeqTCl5BHoH9V3hCNi1u0PrXr1QKNPGjIb
YpWLxRRD4H3QogVfI5BSdmLXdjnelSFZkFNSXGdndNrcGwrhI5Ee/7Nk2pF6p6VD
9kzs0Mq5mK/OD1+Xvlr8FbtHVVDq5cy9Bp44XAeprccgs8xXa+sITHxLnD7Cp1iO
WCS6yvCHWL1StE5PGMLcrXJ+TqU5jUtB5mafAl7Xs+9ts7sPaUhrm0rdAY7zyQpx
GdvJilYiThYzCQe+eC0rN+RQVzSc9i2H/6s5AeGdttP35cDCI/+QbhiHle0iUcZR
hF/4P1gmWq77QEQYnsAhJ3ffZB1hFf/9GXTZzUnwMb2aOJV/Oq3zGVDnZr7ekJGJ
vxe+IP2tnWLnScnAMYmXDcSTFNhtQWQ65bqAlQQwB1MR2lEE2Gu3A3LqZgzLHdax
huFUCyQtzKLht7nEp6/OeZoiFh4uaoLFwtwl4S0b3TU152g0ec6ACrig2YXPIjX2
1gmq2TNXOHyu0BkDcLVWKABqWWcTCJyUCDcjNAns6RiC+49QVs2pS3p7jt/jKXd5
z3ywIoYgj7k5Ntm3jL5hvwZtppD76tASKvOvxGoErtBqnn615PSueiYKPKLggh9S
u9Z8P4cDLC1lYBR/3Ems1pCMkW8BDQGgP3eLYH4qldZ7hTSpZIhz2UR1n/ga+gmF
fWPBLHANVKQlnK5eRbD3ZguuC+QfSqUlYHfVXm62hl/Pn+O5bELqp0gyQBxZNJiu
0SSRRT3w3uzma1YjrrD0kudFlLLGoiDRDep6yPONvXxIjLL9L6agKDTXauEv+8hr
GMZXgKauInNfA/HsljoIjPz77qbWYb75x811pzLDHk7pp+tumGVGmEs6rwd5luql
+zYoszkXVGQiS4fharWpy7rtriWK1P5gOmmASlSGSz3nBIpWuU+kNwViFRViKTCN
ro99Fv7lnq/YDwiFIdtTF6Uo5YsyKZD0nfBY5dr3kKAz3Oi9Lg3IhZWLNyTnVL5X
Ba0WOA642Ae0ec9ws9LorLPxgUmL+n0sKFlh8U8y7pwhoGVPgtpJj8z4tNZ6Nwoc
fyZJBrwbFydjlwB5AkYyVqsL+98Qg0QjTyY/7B2YwailDJV61vYoh9adZqXedFLV
oITWM12MO2mTap3HOJ9s+UNQ450LZmywrCRVEsyzhjnF2CTPemZavr4QCoBmUJiU
D7XhT68v5VVlG0l9JxPoNi3t8T8L8oHT/CJDG8pHejhbbbK1I8rc18jFzQnag8cd
AuHQDO3Xgi0p8l+xWJPAPPFuqigeXVNOiQIvZ094zUurCzCvkNu9nyCuFkBZcbcm
IcoNBnbfD504FkUaA+/JVkgJ/M7TilF1W1LFBQsidc//ZBziJpBIyziEut4G1iTg
tApMxJvNBuL7DanrxRhtJakrtJfVziirKwc5T/i8sGYgcQcQqfuR18Tg082T7nmq
haZw7pWzV3bRoNN2bzhm4yHSTDjpt8RNdiBm8Vmr+PV7ENyo4ecLPQiWD3Dh5D4+
cRilByI9OZdxutrKTI5DAOSAJsYrrkaLKO/Ejk4VcFmQsdGOrwdY/W7UPt/+fXlS
2Vy6PzuO5g58yDyMs8FR6LudSvv1FEaN3dIA6igM548K6uYfGHJmAWvrXcpQx99a
Ci1w7XnWyPee5hRatMqrTG7IWv+I6vrHUH2V0H11BL8QZCNvVMeq/hTx4V5TXlir
YXHI+yIIDdTHYYCFbk+qiQwt07JDCou1oANOiVt2VWnKbmkrOiFi/cRjs4+pFb9y
zKAAguycnVFsv+aBFSSGKg==
`pragma protect end_protected
