// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HMBFSfgVRo/8wfof9H6BW7u4bPziclScQoL4A+N0FW3WgwlLKJ+0KIZYGgrswg4mHa/u+luzhQWH
doZrNOwsnEj8R51kkekDxlaSBWP0//9sLW8Gag03GxbF80igCw7QJUHvZIaNeVhu9eLfZ+7eJJPf
GRyxA6IvtbRSHVOetGD//6p9wBf+TkpXEJM108EobwALuwSa4GLSWLMTNYZhAULBUzv/6dmNdlkC
j/1yigr4y+HGQ/kBTkhAK9x3V27psM9+EGb0Vd0q7mE88XUX/I55EC/7MrP7RN6QXAE4Ezhx673o
LnyHzNiOHivPGFE52yLSjYQwMa15gX+xFlw1gQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
PRUPumx7byliguXtaPra/5Tv6JBDwKvh5gzygtV4GZN9b32eIxdhmXWkYGx3+3wfIWUSy/mA4LFQ
AiJLgIwSDRyOBqaPaHP/83YXGf/YTRlepBWKGWNYe79N/aXt2qUb6TPqlHsH0qvzaQjGRDuCMY3C
ixKO7hwiaRuJJyFKhVwgheSuU7mEAIzhhfq5UwZwms7vz+JC4GEtJ1kJK10dKr7mrPEEPxWvbN/o
/6NdpFn3o2+4HLKmjhPVtPnKX78JaEcS4NNR+kNCUe7xKd3q4hM4tBLMosFHmYPS1rDxvwg7ENvx
ou4mpr2TeYez5A9+9pjmHNE88Vv09gPX8cF2Z6ResUSQ1iv3kDSax1mtUwIp9n5RhhbkVKxJQK0+
Dfom9C0FEII4nZDiKFKrXDz2ard86TGBSeXeyScf2dQKBFKkPIXC/nFH83EPD7R96758yBvIcLh+
leOub7IWMqbyJKtGGYu4kg+sYh6U9+H2yMXh6adMRLqlswRZMDjet+KLWrIwYp2/luRvt19dEqTS
gOzhFpQCg5ufoYzGeIGuP+Uae598nQbvRlVFXMbfMluTYAhooDAq8wflDhgqXXhu0LbixSHxSZWp
AqmXH40QaULXoKRFPiyAJ8W9ITkS5PM+l6Vp3+CiU/DWSKBQH3ZlXMEHLjI/dB7jt9fleFl26E4Z
zmaSBAOlvAECIk5f9GDgYpGNx9zhrJxcaDOQsPZv2xp6Tprs86TuR786n45cbNXjIkejz5XcQf04
0nDWDwLKcyFzq2s8V+LeVbqhvPLqnMHCpafORLAtbPDbHEYmK9PrDkZfB3cOWt6liuZWkgSdNRQa
WNZ4a+KeXpSBo4sYw5LDdaQrYiiGySncRFv5lLtLyTz3ixaUjT1dephrQu6VvPIArFr4h20nSgFh
Xr9aRzwMOhxUJqAyFXe8fVYTN5+wrPBR/b9Wht1ZzmFNMfnoLGv94DK+li+tw/V1S/afIXfevBg+
DZk8CnzEjmzjeBEVlxwQXLFTviirv3d2VRX1Eq43kTpu2YXvjiYDOdt81WT/UEOjlgEoJ26YXMGi
X0DMmFbfMQ9X9vAnnBIG70MFx7XdNO6QogyjODGrfZH7FMvdqYWWKXOiB33A+U5t9OqeQKPs000V
sWnyn3u6Qs76Odz+I0BNsnE8hTlfoUcnXwnHWMZtURp6T8Bz29hK7L9WC0bSSmOAcXbRc39SWnAo
0YZCbiV5FXGdPuZZUV8Dflsd5EOnQmccU9rVH0NK0DTHA9kjaKIh8A7hDqTF9Wyo7+y0cZXRs9jz
qffHcdkypzAmc4xd436xukGEPPH5yykYIqoxXpuFzbHh5QcTQDQ34kOYDGOO8eQwSwrqdMMMRfgx
iKtYOHgo9bqI8TPU23mJQiCobRdE+JfA+I97kGIQrE5BUQXiF216FDTnj40825or8+2KoZzBN6x2
bCwJHUCBGYcYjD7y0cdT2AmBwETN8cgYEX4vf9agVA7AiAuZwR3NIqdv+0Q5I37oQvAX/ywm6GAb
ojxYrh3jWz/K3Q3lVjFza/7csb3erl1tLsu1KRFs8EmuHCWo61A8bw/T+o4p7iUsLSZ48KGauDMu
0ovVUijDIbDUfvaKsXdPWmZnJRg6oPfsbpMEWkx8FcWfoQ/C+MipWt6C40amGj3ogYRhqvBFpFEs
ExkGr2iHQ08Ac9eraRrpsFpeWpqvxDGxySELP1TMEsqVrgs9hUSJHZOOMCBshL6DMIPQvENoF23y
kjHkHw81VSmB1Ea+BF/B02fDO2qL/C+XqaixeZQVWQ3zKHSW35QOCB7oL19slnCj8+mQU8/Oq8Ca
ZnMxYfO4ht6faAJoaFo5HhEOBDnYtOT1d9FXE7AFj51HGgv18VOvWZYczX/0uJa3rs+NZpZFQc4i
bl2+tbO/YG3z/eMkC8FWyv6gUvuMshIKRK81mu/TTX7AurynZKsoaT+pV9BCVIyGXzrej4lz1F6q
tP88qpvkEtvQwQanRr6p0Qg4ophoGeUKgO4aOkFuksT/fUJxRPY1FoVxg9j+WGkaRD9Lpl0XW467
w8RtIrcP4JSet8Ker3Bfp5AhfMxcifu7ZDr2O8UIcD0PYtu6mJVzr8t/b/Ssj1FqUZC0Hne5/gyf
mikBSeekVCvKggwlcdVrYFYjzu8NaotryaSNCO/l7QUVauUejHHYZXt8qyf95tLkwtMIvEAIWBXY
O1oH8VPtouN+ZQsd7PCtbebWNGfKBYU3xxCj7OOmScyuoHlN7wKnXL1C9cuthnoMBnOLStKrG3qP
spuvC7SECprnB3tMypF1H7+Bvbb9q6y8La6RJhUSWtcGteNtmBCGU6q2lVYHZjDZ4xqMnwpy4ckq
In1e3cM8o4sHAioEAN2ErSb8Pvb944lBG3gUN+OLvU7G93uqRc7H2Yx04ou/4tmyi4zCuBcpDR/y
ku1DR0dSrS9LuI3hIAgMbhmJc7/Tfe8lYeCe+g1kw/PS7ZvlIeaWdzK5//KHjix4keKNVBFt7KDs
WZieu7YpK5XFtbsaT8LGCt3uFK2AzTd8+ZXaaYw2e7l0dNvIyuLnX+5p9Tq17nD4Qj5EYZUl0RD2
qLKuEbZqRT0Wy7ajwbSnpclvWg69cT3Mc6U2W5KwL7vjsZZPWcCJ3J3CRPD0/XTnAJWRbTyny+if
HE2dELFAcUgb9FUW3LFTqFeoIPzqwI/Z5bafvMoTeejXdxbwjlkNayKyYIdEn96TPkPRwtQ+xiUq
Xng/j7AxTpS2cmaJSbYDhElX6nBN7jTUy1W+Po54t9iaXle1jMYhii5KYCKk3MwnCBZ3sZTqlTvX
seiatKuc7g7RYIvLEVETDZLJN1/8rLdo2A4dhdqXt5f8rx0q297NDWvDjNOajAbahpN+V+FjTCnG
cQ+iZOIh23rZfBFpFXK6N0Jrfn6k0sI9KEO/crypLN1Kxw44lSYgN0lceSjvdv8Hh5r4+ZU/Ws/h
9sbsNKvia7FJwCRXsioBCBkDj8+w9aDLsH7A0fIFreYk7lE/CRqjyTCXCc5bNmbguT5mh/QPsO7J
p4a6ia/geKzacbUK+2TRXFZdwhN68Haxf/LyUe+C6rja160wWf5YWS7eP45Df7d4zpI9dDUgSTVV
4oLScrRxVcniBE+LXdpH4rP+sDp3NzgPeSOhWMUm17xdoN7pjygFSI3ZZ5TANb2vsLEOFS1iDbRY
tlvbQefeOxPkowPaZp/gsb/AnnZGlcjfJPZUf1Ascue+qu6FlmcSCl3HgSS8HrcuRfVhaD5KWzaW
TiklqiZbB5ZvU5CkL3QRpN2kQ46/cm77dU8LihigISEvWF01J/xjcTePxpunYVo3uh6lxUJwaHD9
7GOVVQsqFRtZ/FLI/CubbtQf9kEPra7Br5vpmwAiUvxCbxdzvQ8r2gJ5BgnlzgSXeDCMAaqgOIl+
quH9xGVNpHwBH2kGqbjGaipiJV4T0inUNqQcvF5b11b8PUOKqYFk/HeAqnH7P2Kt6IhXNUUmxVda
0ihHQk3xFc2+Mgzqk1/wDmVPalHnisSBfRcLv3/8a6BkZjAfJvPuLCYJ61DtmD+K+yllJfwFIFeq
D6WSYvB/U7NKhTTtg7fIXJGPi4mZdTYL+K3+xLFkXtatHsRWAsAFGkBqcxYIdwklOn4lMxBI36zh
qRFxV0GAlM4wQNyy2MOwb/Q/eTnkd9tXsY035i5+iDAkj0/bRdJGNQV3awEnmhqjxU0G/HSX48km
lCRaivI/o8u2gMRm6IWKblJB2471d/NpelZFTACUddENb0DgCJVEDvFLQ631LmDPURAEHzZZjOKz
iyWzk9MvERIPXB1GNpryyzR3r1dqAIIlZN23nECDKq5lYjaQz/HHyg7aDYYvJOkKkF2NehME5sdH
3O/6w/g4eVm8qnRVMpptfdBXkUBecarXVcsDfuM5S4W+4LU13wHTd7N/zMSo4J1YgS50xFzonaI9
eJYZgRClrNYLkggunFWcf5ocdP139yhx3GcXXaSVpkiNKL0CElXJOwtBk/2ONRNPjMhhPOQiwZH4
OETyxTKN4sC+qqvG7zhO2NJhhdVUx4y/P/RScVR2mjQL5sYeNNAoqyF9bvXsKf613OfLb7rsL8Yt
35qVJ6VTePYVL/QaP3s6hVB217qwJnFu7aYnSFqFMTbBFv8ZmOWmnln+IVT6KDMeYjJgb9jY8yVl
vPzbZAXItWscpVKOPH52R5YsGhgzsphJRDJT1z9x8TXWYPC3/Gr0RBLG+Z7Ww9DDC/gwh3UZGTii
6c60Q7Yu8QQHiERZJTGUsT1ZFFrchnXZGGYkHaXx0GrSgWi9EKuuT69lNpXTZw2NCg0Chj1bjRMr
6IAIWYW1WywKHjS9N5Wa9olm99mnQ2Xlri2VWKmE7CWUFmzVhi+TWRT5ZAjPRS7k5U/GtKsPkPk+
GNQzZsA3eOf5msy+NT8ITz0InNE8r8ijw3bw+SePVZTKv5jBqEWwWSk/5vEYyD6sWTaeodBrsrhB
k+eX3Xw3F66W4n6Q5+uniZNU8helz/9l0HtywEjkGQFU6quDRK7Dl5kQ9yzGhkMsT6LX4tbKnive
BO7L2pATRtuX8Gm7wIuF1iljsCg9kwNK4SgfDRHb6yocdGu/HQgbre+uxhqBmdLauvjjseZfNW6J
N/rF1m/480C5Pf6j/i+t2PCQ5mKviqQe64b+mSSZqhyoApQR5RV6qSjjqpdPJl2Sq5/+1BRFGKju
OyFoUuT3FgfREDZ1esr++T34LCCdMJ1u8nVAzw2REoqlW9hA7A3WeNpoPNL4Eh64kBlbnXI6lQ88
43c9HqDfFpT9WegoD1exvgIvWvzNgiwZ5Yubn4rMaLXDpXlBQmXttDNU2oqAGJdsaC6HVRel8gBQ
lpTzNeHMAyPyTRfwYVYGKxrBJYyzasPNP9jiI1gY2pguq6W9Ce6niPgKjgyBr5RDwlCIDG7Fd18U
o1UcBYcNH1FYH2vvml9Ie0/AqDI5Mx8S8fX5l13BQQvZTDiRBlaA3FaH0UfzA8KrlR2poA7Hur+X
btgT6eZSHwWzS81rvObhMPoAj6wl5g7tt8Pqu/NBFqbTbWjXmh+5a5vNMAKP8JUFWOrYIEWQkwf4
GeTNHOKnEsRKm3UGUPXicT694+ZlaFwOAI4nD56w9yIW/fgzpu9RyU8/4ZSu/QflW7AqNqUOxGls
Q3dGHWygyvRB1sUoXuTmNrS6Cm39uMkJMTrI7zExaxCD+F6hmF0pK1acXlTZmRv5VoH2X7aoVNvu
YDEmfKQXLQgSC0aLJRzpfkTYC/vo5Mnh+kt3BaPqPutfQ9S+DIAz6CAopU5k5wTihrKcDhR3EU0w
66r8O2WUKnw/l1JMf+ZaOEQU4v4ekc0hqvOuhi+CJ1RTFKhtubhk8/GvRPSXbs8aEgGcMhKu76Qh
rUkHa1ELkAtQUeTrevR6eTGUT8EAjWJFHaf+/jFg21RQqGu9wezncJB/bbCHTuQ2mig/0aCyAZKW
BEE4C+z3GuX3ZedQiMX/kC+fO8RIMXHRYk8/Bvg+tBCE9DdIlUGvqZ48pvyK+maMswAwffUJ1Zp1
71f3fobppGV2ZPS+N5ymsWD3qBYndhbexdXFPrS1kB/ZbM4A70Q6PAJBT7LxkHjXiDBSKJ+eSbeH
jk1zGUqLXHzyi9u4+gMgf3hLf2FJ5pXGAqYRJurBjDF2UlEysPIGE+Cog6P1Do3nuScDJmT+TPIK
UMpZDW4/BHYZ+BBXQsGll91Ae6vnVaaECL7A+/PsEl5DLyGaOCXQbXquudJtnz3Lo0GQ/0UzGGy4
6VuklmZxffMCFDV+ry9/FKMjxRLOjyYBMR0Ppy1zNkMBCRTDideO2/8WQbKpKGmeUI4fS5ilXmdk
lirsd+YCIyzsSv6joabOt6qZUPP/902wAWHczsmqCObJRNVzKJiBNsexGfzMrZExolyt2qwoxHUe
EaVREc6H8oQohYRcErM3PcvcQsP3qXvzHwNs+OYc5jaZ1HVLAera88DRAAJMsXNAq20uaozP/51C
kuqY/V09MobmH2foOgBpcqNOY+VuPvvSR4UH/+dwfi4KJ2uc6LSnqRqmX5d2gOBbYgr7C/kRsin0
Rkhl4oCn9h/X2usIQHQ4nflzH9g79oKI058pJPD67pgdSCjsiBAtcJmXCpNxEfmlEwrlBx+Sgiks
6WWz4wZe6n5KV8QSx/gIhJ3OwxADn9WEC7LTncZ5F4VngdAeNu590fiUMIJ5Wbd8oQzQYNkYnoyd
XcN9O4Ei9cRGlz/ESyYpBV4rpqga7S7oQ/lMr2P8spYtePSonBFVzS0THlPhSYCk1cWf4BXejGFw
OvDqIV8BG/TLOgXkkPkmB10DsWJlvtAJ6ioHwPmgocBqckM4YeaxG4GHzhh0z2ET+Mx5rIEKNy02
2/M/9L3k2GkVsMUXhRNkFiwrxNe4gKAYHaBF1HRGIlLuP1omKgCnagTAf169Ci5E1CWJDNGhkHHx
Qeg8l8kLYySFMNL/BVdgz9RGHO2XP9Irclzf8ko9tMyVpIaZl6WFga3Ty3nxvShPp06arkPpzP3f
kyN4bUYbAmryTz0k7wCYll+vhJsxhdp9TY+79O6xvX23zneVvEHm0GvnYmygcOFN7PzSoO2Dv9sL
dpy8lqavH4vuggFVVq1Qy5+PaOWM471FaobSdqvfi0betEdIYC4mt8npMB0MwkwSf7uTT4lU4b6J
XcxBFs5CybbVTKMcYEjGXGQzkgkzrGTjPSK6ujwAZL3kmq0D417mRelEzuI7v4O23W86IFQhiOdT
43Vdkkg1S15SVeEK2tuGIzdAxDmaJyLmS+sOzx1uxnV2TVCC2OqgwaLZJxg96gWmuCVi43a3+9kA
3+zuLITfkyiFYZdm2wS7MX0DgGH2O/u3piGmklRMGCyiJ8+8w2rPO4XGaPNzg1xLsigqHadTKmGE
IKVTPZfHcPNqdjmUTvMJ6C37UOFwtCicpvtf7ZyyCpoJppa8LDKi/tJ0R1j14LMWCrq8LN1b7UKn
PXk5fcMHwjkicmdzYCiW76ORqrdmHOnbdpn++vs+EXpzGIFZ885/coS4biVyo5zjBKHFpIjlSGGM
kc73dpeTIB+9R5+ER0ZGNkzhREKGVmwJpm5JE1ybY6NhBQi4ELbnW4rGfe4MmLAJXmWi45HRrOHl
A4AJxDmaNh1lUthhCP5aZjBnjQ8zZhB/+w1zIXPdgCYtnJb/5rmFt06R9EJXGju852Mj+4gNlo4Y
MBaaOh+aQ5ffviAOXnXoxP2lAs8g4HF1Svom1ztDUaREzRzN3RxC+BepWoZ/ZVxAfXjHEWzd38XS
FYnG/1pVRuFvuHg/Z5VNdSTb9S2KDUR5hI6WLCUkFACfiy60S0WzrH4L0f2hup/AvXa5Ij5L2RG+
1MMkuJB3TPECKWiiCgoi2WH7gPrdtQgBIt48d7i9daIMuPecv9jDeXzkAesD9Hy2zcuyDrhpVG+L
yqYDh79mLPMDXB71pdLPhEf+ZzcBe4HUY4pQPzp8of+PNk2gLK/poNwaiJQSGTdwMNMQCl0yCtf2
jksDuaJS7FKMPIAsp64dFU6ZFJ44UkbdDYcW9GcmPAMrmAxwVPnKWH9mYQJzjS2/GQrqN2kVqXvB
xFeXvHglXT8WtYX25GmqvO92RlwWHvYe4tQ9fS/BsD+qhn1/mYXKl+QEwsPlpWm+4BoSseNulS6l
qBtDk87zsv7RKw25tvTB+9AO4Jz7SLnRrbQaOETjVptd/nd0czDPxYB+7gZB63qsyFlk0vdDd6eJ
vbRLDNbAnOddzrfTcs87BbY8SkSdH9n7RKxnpEddbVqt/FkPwzcggvm+AIkpqr0wnJ7EZFKQ95hE
D05+yRaOvXEdB8qQjrHdLCUIG8CSFXJmhiwQ560AqVvhAE7WBfEfH0CAsvw34sCg1IPQ0qSfcny2
jzbsd8j2Xc4aMqNrotEq6TMCcCgtNVNfjZbbL+UPd2/YPALB2MFh6gkYrimvZhQZfKGP8r6VG8Ul
HWVZuH9H72HMZ218FJLdl4Aw4X1VRGctKTBT2y/pHR566LqGH4b4O3NDPniqsBNazjAe0qoWWMq7
k8nDA8T9LGjSPjhECa3+ZQDtY9GRf60BJ0ujfQ1gSiGK0T4dynIN4t9DSIeCdO5g0P9qAHA4+pBu
4CP1V83mYjb1y0mLrH4aI+wxq/lg6o+K8ImUvq4YBc/8eTZXxTOGg0R+/s32IPmLpuml00DmXuq6
Z5VBQzKEvIVInILMfmb+UTWX/7Jq7AhNO7PEwO1pDGQn0vGTYoBPJmYAxfCEOgJivoMuySgCWRm3
Pru9ZstIHZ7IHmFEMUMeK3V3Bfzv7vHQXExp1nmFIAto/EEQP5+C71SxkzCYmUz3qiHsFVG4LHsa
+ceBawayM5gHvgPs4A5JVTObdchqWK/gv9yfOOQSuVqAhRPPCH/jX0EClLJH6ANtAxiMK7exeRXB
s12WvnItl+0XhNA+sEZfu52kObcJp+9sTZVDbJVHAcO6s3cJfaXQWR5ufxItAKonKljoNEmYM/Ol
pnYL29it6F7YeeavJKYxN2LIDP2H78i7OC2t5pvS2SqMpVTnK6SHZ63ak8b+acL0Hn9UTpDKlYID
UlwlriMqrqEw9OLjYdre0GePb7H8HGdpEH9x2SkXmcxOggn5qDlviG1QVOUUacn86hBJH+2swMc1
qtFkvn280tfGtsAmEmPe/lXistLUyUAe1NwtqotFbWhoZDyEpBV3+LZy8sFYOH1TU506l/Yf5vKK
uWpiD4BmxahpBNFpVFOUKpMvDO/JNzBn61Rzwtg8Plulx93NMjrW+YWO8e8LQGYQgEtbmLLSioqc
B3IIsMeaTk16P5LXw+p8pSF6hJdh8qAW6F+laKx/P4n8RGPpyiqS7Lcm2De/Y9NB8I7ILhSgOI6u
mFiHx5zZfqaPMzUh1WXLP76qLDePO6huVpDxbzgJ1Fh6NgeyVuC4ZU3l4dVL/+4HH1+l1Bsm7EBv
VDhR2qHBq6CknNzpN1HT3jPQpoZGEI1ImJ4IEIYJMAqAKRw0HFF0+CsAPyDvMfvQYAyXoU+pExzb
mO871kR1+NaeRva6mvIxaaMlK6+1n9hDd8ILPsJXZYiPNJYcGrzhSfAAtvJJWh9JCj8yKacbjLMW
QWvDyPuMxzVxN+cBH0Y+6ehXdU9LfsMKYujMHPj6gMVMfnuQkgaNCRPDRzOpyImyfrgYgt03QC/v
fTSk9YG76KySxSEpHYmODh+dCZdRRNZQen1dkWJsW4sMdXnRCSRhG7EFWNu4C5A4Sos4tMOOd6m6
Uq8A6dyoPFAl5RIrhmhanJmUCE3ea5RCmOBbqIUcYG36ulc3RnWPh7bhXhgYG4ybh0ZZ60pA1U4a
u9jVEIXw2QdXqgNIoFrlPkVR5HSsamw22wD8ONcvIAjTzD5REsu63UpgIzWEPk9IBelfg48E2dJA
wR8XelfIAdUWhJav3clb/pp6ul/xttgwUY7CdV/H1hjBEp7PiuG4IXoELRjea3pmcBgyht4n64fV
qZfto/zDHgsdjr9QKysP4o7p8ZcjO52/c3Yqsr9MFlca4zGM5hIvDLe/G9dg5EYJou3j28FITEr/
uMHMGyEQBOwr3V4mF6hFNueXdkFzvxoOdMEbMLvU+s6qACEZLP7icFWFKeHMicaYQvCVmd2vPAXG
pIHk2bEILPq2+lu0mamVtprfdSu6YIteHzU6wKr0G6+qlYg08SHZ78qD1mmRER1H3IAfR9xaM3s9
zrOBEpS5C1is1/6a1JMT9cp+epJhj53ZbRBEvd/th32RYhErYIl32UK2iXtLt3XRY121vJXLRgCz
VNgmw9jz42bT5XE0BaakFstAjzKDMT6Pci2fQPXs5Iq9DqrMHDEHjvxlTJKk0rzfdMrchxNgj+3L
qmC1FbqNWN6pXV0dpcOtA7Rsob6s9i9camONmZW6w9G6ItJRjcF3KyfzgFV5yRSmKKksFCSaX9QO
qqkwlGQfcj65WVafVknXdau+TI7vpH6ywVSc9LN25/TXjxEjvcG7z6YjHKFd5iGOIn06SfW1CNmU
696+RTyioCHmKjgAlqELY6Jrmu87goVwVJwF+iAFadwe3P7VMYIWyQgzVb0s/euDdnRMn90l8R9s
DRGq3rUxegaPdLfeAyE5T0epEhHaoeIoUdEKS4DebNQfnl25QsE5OGWTNBc8mRQok64ATMtU2bHT
ig8mGI47JKA00U0vqoogYXRZNv/hwK5QwfwYzNNSxG0o2vmQUPiCaSS4EI8SQJzgB2zJKMxePV2v
yKncC7zZSYYnV3t7sbLrlhJhSltTDtl+asEfttR+k3UEfQe/LBiS7CIMzY0OKk2ibETJs7p0mxX9
ki4tlWPZIUqKTtHgVkn0cp1T28tqUS0RsdPZdTHjdfcv9ub1sWwy7fuTwDpp3gydqPKfNf38bIFn
sTtU6WYQPxMhSjGzuMKfVK2fC2f2M8Gbf5TFMELIDDiie2khKlwl5AcQ7z+/L/7Ig5KgC6y58Jus
qE+a9EFqPPFDMiI56B2NzJA5Tri8NkTciMri3nNRoyABaBu+GMM+rUKv8OPpQBAvV5v/KliwCDXb
mIcjEVWh7+3mR0je/R5ObH0E90S5l/mPrWFyHNV4F6fV2jFBVf+Xr8TIMbQMF+B1HBugpelJh/qQ
3I7wbmDoMjzhf9+UpCR6F69MX4AmtC58bxkYsLQ9qFkklGmXRiMKdX8fuBDUg8/E1Thhhmr+HIH7
Ya2uZroDjA8IoO8DmbIz5wY+TMzXfW8ABghTH+ltL4ulf8w6YDsV580TKgmDYebYuqLllhJZeR+4
Oheva/KHvdY+C5z+I5MXp6XqOO854qublsX94PsXVmJKGGXTmcXToKT/qo8W+Kk2tzo6Nz2r8G2b
FK3+FRcx+dAMCSQEiU62mG+0cxSBUogYQFuZAOOyAL3kRchWrWgEhzpHLtw6POQtuLcd2ELGB/lE
MVc6cx3wLuKjYQAt/xJxfdcYoUWwsWkGb7JrF4O7YdTBkSfWjfgH1qYXl91F/pfXKmPn4GP4Ukrm
TSNTGpjuEWR8Pjx97KWTUeO98npCrCspQJosuPRZJPhCV6wnIk1KRSy317iIatGiMYmOqOuTybt2
XO0iveQIFyI945chJgBDWCEEwth83tYWnY3sYEhvKIr8PE63K12C6czOD3sDDjmbum4zjS1xKtJM
xclMMiTApc1ZZ76gZ860vCAGt5+Gru44rzRABiHS2Me2lk4oyokVQOkE8TYzBXQ75dA/wfdD7MFY
cfBfEVqO6sc13jXhn06KqhMYJ31rXFmP8LNyLpFhO/cb4brmUC3Eu3zN3Qyy9Ogpp+pWyk1LlA/v
vcveqpBPSSotqCww1qVYKZof4dGGFkNap/PTGqyPZDpTv2wxBzdiEt/yrfnMSzTUzJ4aTt+PjVjY
aNgR+CAC7iuR31HZ8DFQTXMOIE1sy3+e4Q1RTLsvTtXv/bHhJ10Njzwh7c2DCre9N0gElkz3+kry
ChX+Fi2ymwrI8zW/jiOM1LlJPBTCCaMO8ap346lsWlgCx3qkPHc/LbyHHLF4PxaienwJZX38bs+u
8MAkK/cqFy3EPS7mWrmTRqr/rbZ+sUfYKkF3LXV5DJpjaqy+7hT7hTy9m7MBP/iUlneF4BiauhjI
AbRivJJeKnfQMNDjKrpVumARDK65bMH2Z57i2fTe6v6yAtimKkIoQ+ZhoeXjkQM2HVOBnUZ2IRdb
uVUIWxN+acPP4pyxv8VnWas7JVGZPDBZSEqCtSy3BjIlw2Z8rGB+wkJC4h/E8QxsE7DS4XBi1COD
rPEv0ZC6QweTMDBwN4d0hOCBny5TO8UDDwMMCpHZptuTuTOi+RI+MpFYdPipbmy446Gt9Y2IIwtx
3GEtNMuLXNZWjZsnKKzIvxGCz4VzEHQ7DsDNcOQjUy5eJ1lHpj0gmQ28223Yzwta3siVVvyiZLen
wMOmtkijnPSoXLm5MQONeRWd3/NHBIPwORHVtGqG8g9SdIeVrlfjpGnG0p4zFLLgrCLw7nRlT2Xf
xyBhGAAcfv2mIkkcsMQMKdjFTD9QunoVDuKE7ToFrNcZ5WCux1DEkepSmApXu62nVly5IZr3d63y
rkniVq/pgTeGHhdxDvfqiyA/W7nEC+ku3bLvo/t0oxid1RJ744Q5bS6GVCKFVljdRNLhYw+5E1h/
k0tbH01f+kby9utqGZnAdTuA93S2SXdbL1772Z7cU3gspwD3jjITeeHG8+Vd3EY3zwGlbs7bT0om
rxZCRijFwymWmfFcD1XC+tYG+Ntsop3vNSP2vwvRRhCc5VQ9+n1gYyJX6Mt9YFz0gl9ReTsx+D3T
IhdS9YApi97Gmyo9qEks4Vw8mu51/2WEVrXTZC+JVdlRHUeEZ0XVFgebz8W1hQQflRFDVhW/Hg2U
+JTkIpEGMo9pk0aaEAehz5Am1SFGFe1qurB6SnQ7/qAC9wYBc7biI52Wh6Q4iPm2zjsen+7d9Nfn
tW6uIEHW6RQDA0VTPmBBzzaNrUKacIxg8eM4SS9M1lPpg94SlqPFa4I7ww6n09JW+EwKQ72chv54
4H2ydpdW/o9mDLmv2V+fSJKh1D8PBG02GLoC8jGO2RRiLGlbBYnbriSr0olLtJE93K/KtEGPEZ22
WWXV7g0/pG9uXfuyftGccVIgOIUoaVIYu0baQZNvWX0YtNuEkJlshYZrpmwW/L3owuWL1oba+Xky
/+Nu/JtsUmDll3FxnIjCLY55Pf6bmHpalpwuTBYzJE17gHkeGXP1LDVeR6GmlgunqROy6GWAjgYu
EgyZGcn8zN8kjruhijQl3hqMT/60DaQ/0A7aHpJeD+AKbW2cgi931ELAL8OG0xH0j0t8/Zd+Vedz
OvgEY4QSXokB7cjnv/0N74ZXF97dW4lsr3tCUl9nizXHf6zAs+jvcd2ETb1h4VWgcayt+7Tzleft
rgDqXPFogmdQXJgPozWXf9nL7Qqu3S7uyccjWyhYVMlOFljLemxA29F29NfDuCG0dQug5cjZam86
Qr1R/F4vzNRqlPxhaDATWLOkiSHvOODBT4HzfxiKuWnmmzsj/+rTIkHKuotQkZ2g7UjfbG87V2ba
ovMA8sJwX7EWuvpBbwNjytOWxfBigc2jO1A0fJcS7lMvoKrt3zbUW/BwnCVLW6al0TnpxBV3G9Ed
SFxcIKESvPQNGOf41J+8T+t9deRS6/I5R/COvx23vtP0i6h2xCrXRcXDwAwNK/xZODL/NDWo10Kq
PT/0VN60h2MShrXB8qByHCUxv9bnQGopm7p91GMN5krVNUI4HhAkSl3zLfoSVoVZJOJeY83L3tmc
UQGxe1LeIi5Mqa+I1lXjajGDRO5w5BFEBtAxojyrOttQiDQDehqSla9veQ7hj/FxdZN+7F/SlhGJ
cPQACrHT6fa3jk0oNTR5ty5dBuX/9Ac7/SY43+75QVI+kIby9rzNDibFXn6DL2X3NMwogzVEmu/5
3FKZ/fNbnQz5m2m2Z/WBnaRKMwMvEu3kM6VZXcW6AJ83bKZiTyZNL+LiozOCstOE61RgQRVGYrSR
Cz4TWk9kHY3bO1RVkhE9deObV+Rm6rus0liaXd3ToTUSSY81MosZM0N4OAFVrXF4b7lxG2/xRicy
BMFTQCDtp54KBO7IvDSVDQS0rWOFicGx5dTYKYcAzotNe1Y3yJM7xqvjjB/WYgz3sJI3DaMMKlUC
aqntXILO2CUiqJWQvbG5E92D0FXf+lNXCkVDIdLEPuSpSYDIes2QjZa6d0MbypyFhS8HDdt750jJ
/2YzGsmigEkM4OYOB+vp2VRzqBd1MaViHyW5lsNH1ySRL+JrL58vcMa6UBTOYlCfWs3aJ2Ff+Ruf
HNAZpobunDpoFtmbay4lW2JRTLGEGF93O2gQDWkJcDoNQhIk7bVnsO5vcgpuOE+oEKV3kRSD8Czz
JVqZ+FvhdGc3SPtisBB9A+vl1ia5s+tuSubIGYeNxAO4CgbrOHaC+rtsmFl/KSYikQTarbBb9k3+
BRdbkafSdOiiR8g2cgaB3ME5I1RCEMOsu6BOzdpIfuiwAVv4qPq47ywuhLoVyIefBhEELac13Wrf
N/TXfkNmDQXhoa+2Kk1TlPGEKQXUWQWX87TpkrJrutC105s3AOuSkcUspsWJtXFFZYMRTU2nJx6Q
RqfwAUm0FukMOekUQd7qeQYIoPqA/CxXqzlfpL2M/nVBEDenvEPuNsK3OaF6Q7hY4KLp963jHfFZ
3AdwYi7t8yCVeS1fPMy0vrCOyakN6If4qthvf6dbPg5LvV9TBaQpc1sYVxpLijGyKkCyfom8hj2O
GQ14USQOs7/iJXM184v+E27V2cM+JLDn1dixEsG1yUztvqNSAmFudcMPeDpnNREfR6L70NBsyUBI
RczpPgDOAgUcbORJ5MW3IqCEa7VApE0OQo9swbSG4CNyUUfgx7ugSUUpBmICaFC6XzIC7ujYSNh0
iPnUEUjsmgVdg1J1oFVBiZvVNdyiLUJKgPLmJ3hAnmpeYvaRTVNXE0E8TKBqo/K/GQDuZTkXeBX0
4kD3ySBsH+B/a+V+XPY8fB6sgjPihSv5+5hiNdyVgXrj1lgE7R80cyfg3I8jvKlABjgZZV9ZyC0q
utri2G9oV7TAtRfQ4pPEf/0oiXrLP9Wc07rbFC6VwaUJYDFeadniTSEeKwBaIYdfNdG3Y68qVLYW
pmqqZ4PG1lipF8D4tnULi/oP8RPOrnLf5QFg7XMWuAK9Nm3nhuXWzd/Q1AZMWmTDpgG7WfKpuozd
ZKFsb0N3BUcx/xlp5ht+jkf1hjlueA4cSDQU08JM8hdoQeB97waPnfKVvKpClCblTUAVhx/MMqqJ
HvXnq6uFgtJQszwIQHdoCgRoWFrDY6viXSLL/8gUNgT7Pavu5WwTySKN6WLhj3wUG2z31Szyufhy
XBiUHahxFLAcABt77qtVEvZc8sb9/iDC4qyuyEU0vHJADLY2Lzc+LCwMPgXSjCvbmLqDSaowH8+H
ubkKZDpLVqGUQ73j1DvREQeKfnBDB3OgfBQciLt3TA+3J86Q527gViP6SBxH0qVq4JxH7/l3jA3/
j+quvG+eAhR2OOQlef/7GUiSkXFGv16SNvb1nEtSzLViNIh35isjVMDQPvhkrCP29vDWxwFWpVFW
h4oJbK3FqyHTm6JcKuC1DrhFOxeQuKqQM3J21j0aqJfq/LMXRQsEHyohl2ZymB+f5HG+rk4A0BFA
zx5qIj4ThzzFK/WarZoyc2wLtLKrp/Gi6byJOgnT4H5crU+KLTEK/aTIqQUlN2BTwyHc0IpNdTVe
Ie0IWnmJIMsnRUOE/6UtmZ10dhiW5GV9euyRkYbfgQM5v9dF6iLrMVyBPhNkgikbbU8UlzE/zHHd
mqDlsrgg/jy99n3Wzxzpjeb/Kq3g4yt/pvYLRc4PvRmHVIvCvfS5YHk0SvAT5gwD3FiqjcIipFlU
e9Brgf0Gs/saxfOrnZFxIq1hED3efkqauEP+GRQdfGw6AJnlUhI64GHEcO2r4gJduQrI+lmK+60M
D5xV5KQyxpD9xBSFqQB+cZU8St8Ut6ppmGzL3zCT+PI9wQnzicIAPp43GoNgvPrZW474M5Nluit9
gsCMJrZY6r3+dsDV5N5b+6JBIIBoMskK30LqeiKRqE+cCkNXH5pNpyiXLUebSHntaLFJYVAwJe1l
xjBBK9Y7YCsKOknyuGpIxswqT0teX4v0DUeHBCSgBoM61OI2In/Va6mMEmai/WTz4jzIc92O9kDn
s5TB50rEAXuga4jEkHX7XZA9kbxoDUSkCMs3AC5yKFJBoI+uTjpgGUuksVeun4AlkL8bc4TyBkiO
nQQblTXPXzHUWNOxOM3SbWjJ0pkkSfBS5CIoKXMMuDbPKbUcwmIQj7nQcdmLzWhxlWkvH4AzExbf
3PpJ2m41QK8R0o1RCJiD5El8hXW26IvFEhs8GlHisv2xKLcg8yXLETALc2jTC7+AK4razs7Xeo8b
DjtcRNuWNAsE6h1sBcWtPgbcXFjhXIAxHFEn9Lrq0dVWtk93SM44xizwg8Tkq9REBT0LJnE3lyS0
N5d+Hs5s/Bu05k5fuMZFDYdxphkr+P0dTBO2scBd+LzHibjSkYi8R63egMFhQNFr5lSNw/CZbXz7
8jwyFNPaKs97CYtQ2KI6XcwNm1BpV3U5ZUyTRoYmsTtfzeQz1nqCdHRhWpycXzgLooN+D0PBe4iK
zKf37lafcVRlnkloH6DDxEGGnPJH/E8/PNYg1pvoM8It+IAEVGe55E3evnNDMcarcPbjfISRJo9g
s9MoGK+pZ2cuEv8ctcywZ5RaxOU2d+HCOhNJbrCvHIN/1/yDkM/tygRqlARt6apMQgBTJ266LDgh
ZmrrHZ2M6l+AFByN36Iba/MfxXZHWxxNvpG1/X2s/ZgK0Bm5l5Uml568lt1o5LBLb2lcskb0fJsv
3RvPzizczIT56Btuuf4r+fV8MyHqDhAY3Cq1i4UtatZ38NlgiH8XUNa5oRewAmIbFw2WggrWUz3G
EABkTv7tZrhrNBbBN9y3RzsT8ESS2sCZLSTxqhOcYSrR2IPPJWapPOO3TIPpD0o1bMN5Oyg+S4Ys
tY/nIniSXRLAffD0ogUNaTDYHXJa0nbQ9I1jJ5CbolNkoMH1axkeLXPtegFVPidVMhhuxlef688n
UtSrH3W9GT004iOv559jLkGqwXhMhoYHGspvzrL0wkUNTdo77sDxm+nis0VYcCFQKXjen/ihg1B9
X7Vkl6mQtJu8ByOrpLfMZrbXzQW2RGTh5QabR++o2zF5tW+zRerO5fllpZ2a5ojqCgLrgv3NMiSq
pZt4qLdpIvExfymbw9i7huGkBIGMHn9v7vCJeXywVwBD1F56OFNwBuXTvf0E2fuAwdoC348r//BC
Jd3pnbRk5icViDcmCtuzo3FCDAQwMJpn93dD4DnvRlYqBZyUuIRYrNRGD2cExO/UOI95wXwd+PXu
zmlqOS0etut79tg6MR7O+Cc20BVjVVhhh0JLK36p8vxQicQHSxmACfHpTTLIbl+hj5h0Kx4v1Ewq
ka+OCXwykzhZsrmnGvYjmuToHRTeVYOI+g1WSNNg92eMXd4sZcQqHDcZ2NcXjwrGijosTtv7CUMj
+/xYz6kRVBctD3iM3ToZBuohnJbdDYD6pAq2+BxqAWIl8HOKyt0CM0GbGznewb9im8IU/6ZdCZDB
97ORT5vgohEjoG6h3tfYIDc9Vad479hjw6h3F6h7enTFQ2aeNwk9H6RoXZr20XySTaVWpolJ4Qqd
ozHmXvR6vE6NC6W77krmAiuZOmBGUl2097IaPazIbnfH4g40Moawi+b2NpmY6AiHFv1Pl+9WVY+Z
ySST2Du1AWc+MC92iA/l8uoJ/Lev2BVM9dE0UmJzbhq/Yj/cHFxUaF0m4/mkZ1YFiQxaQ3hfSPDp
iwZvL505fTppwWFefKVvXdTptqpnKHza1L3aIj2b0lBDtEN4+g/6D9Zy9vJTMR/9Z1nNx5n14nwK
BYrRaQAC+y8dll/lKOg9HCrVC/aIwUrtee4ovyVYmw/RdYoj47xcYPlahfk8MhfmSTcyNgxS8+lm
quV9thAzgdsTF9xgclmqKlPfyAtrcdJmFzT/9XoV2CoIymmqJsfIs//4kxHI3wAu02OqdDztI+8t
O5IFGwIYNvMepSMzZOBj5aKxLcraE0k9eT+/FZNArjOAkJJjqIGNflTTyi6/yiQj/X9nPKlIGTd+
h30K882suoTwc4kEq5NlgNLTwfxtCKoCgOGvwBAkR+q86Ep2WNVgBQXmhnyj3lUdftgqtrXIG/Ap
7qz24qlrQpknxPKjz2NJASM5HyTuukds1bcm0ZuJtncxCCM4lE7Ef1OD1erlmEr67KTFSXvKIgc3
hOmSXSSenXJRpBupgWqwtFAsgWGkQjUz29fRbsegEa028lgXTftFpaZmwyL1OCZSaIM5GZsTuM1s
0N9B3n3c4uepCqUI+hDjWQyVmKOcdk03qITmdYgnXULftd820wJOWxAlUlauhpEXRJVWzXEnUWWU
TBqzYBu8Tb91mEaNkYLxdJvYb5G15VdK/EC0EYAAVm64Uw+aEl0HazBhKUnvW1IOfLCED31MRb3c
PMBI667xxvhdQv6weqGGCzbOHlXqAYK8mucagrDfearoDVJ77TOdsfiDlLbNm7Aat9uwCjJvM2nw
/kervTLAmgXL79SUgj1ujACvVf0hhr3Ijj8gfwtNlApLcNAZEUROjViJVlfGIJJ7CoetoWuqrYLA
t4w94aCT0LSUzycfjrCeH7X9mmqwPXrd4I7pofz941QIE2/K6Ehp8GoAGTdnMgpVB68UvnvyZuxu
k6f2VeAr5JJCDlUqRnaDM8RMG0tz2w9XySypGubDf6ObaD1AD+bOZoHKfnSqU2DGjtPljH6xiruX
tW1EHYL74mSMa2Sf6EPBoAAlNtQF7acPu/g0oiznHWEAmjwClCvaVctiVi7mTy+2aJtGMgXgueix
OhRbJJoxtlXUP2ChK1kpOn571fVqIbaCLAJcrKZtNK8uMez6YnnoqzGkyZL5Nhi6Ijhk1GURmnl0
IukzaQZdtCbQQOGqyQVAy8gNGqmiXzbfbn9jHCVSLihwEkxdio86QjxpYvriP3wA7bxkQx9QrBzg
Ut7QKNF5Ojt8tagizfWlprv6YEn1wXoKth9AsY4uy/DW/Tjcv6/dAGgBn72acMLxOZuaaZp/HnU1
AID6JIenxcbbD1K5vUJNQECdHJwN9HK+nBpzz66XZyTKqjmL1TrK7wIm+OsFLSLgJsR1AwmCSKbe
ZoLJLScRTN4JzkATgdJDPT/yNcedSR8jy3pDONIDM1XgeI4CE2Mk58j0GkXnoVr0fzLzIQs9HEnF
rj2RZtvn+vt/KtSgROehx6otrV8FblB/SMPO9JRdeHyudSonhFqaN5N2hP0WjdG6XNhEZYznN2De
4qdk/Wbhed9H5Y1VtNha0cdHHmRA7jMbSCK/IEVvflQrNu5ZzO67znkxdt25PT964YWZKtv/8HpV
Ie7EE3AuAOT9ZFBmXaJBOeDLtzEAyQw3kywMp2MwTgGqhPfBGDQ3DYLUoBh1yJdpgn4AMVe205ve
DMMzLGr43V7SbwmQo4p95ARd35AsVDTg8aER61V2e8I7lwZ4S3olVKdUFBQf6t6lzBSaTuYCk4/a
lebAYm+jlIWpXiYA7YJsCrpKT+3QpMH6t8p5l3z/Oit9ATeRmqCHZjFUxK6VifILtizPI+Lcjp+L
dGm3dGB0je5gS/j89E8aDoxxxUW2ZT+sFnBMEq2+PJIIJTcdDdj6K9DKZzK3XAye3GFbzMBahtOB
bVSAPKQkdfLeejQa7mUB8k2ABvXGVwVPqr20u8nLh8Fnn4wE40lSM6n+uZwIQsu+NCqw0/djXqwj
S2HPYvglYCvu9jmMjEWbDhGhrJDX9+U7u6UdRxH7K+WnmiiW/uX9Yj+DYsD0sXSd3Cai3tZnDHuG
xU0sCYNEPt70NRSwrNqLq8CRMHRHKitsLaxirvIJO4NhykUA+LHvYTlmMbPbdbXcaHejYxIZumTe
Mo2TrBmB6qeq+MMnpZblUvWDyVJszSM4MpAX5n0PPMC0fqpcQ42tdXCyuJz+CDLCCUhFMNOmo8ek
y+j4HNDlNDIzyx7AXAlP5NNTVINqsUfRyHjRI4USqyynKuK3d2tzuSratxqXDKl68n4HPx/GFK00
rx1QEisxWn7j5CUapdueKOer0YRNiX/U2bTXdq97e930cuaTCgplpyIDLI1OPShilGd99qtgPp0r
vXMWAzmx0gPZsvVKZ9xEoUWa+FDpcgOW/4a1EEcVjuSpOldQrxorBmW21P6jjOpnPEBpOVTY+YTp
dTC3C6nGBGgPXx/ypYI9QItQHnjXRbyQ5Hl49Ohxh+lDjxSEfWRkBuZweoT63rp5Y8lJhDzlFX0P
LGJ9zA3Tr5NoFmoMYRw3SfqmrbiPytn5ERJYfiMVTh6mCVP3Od3Jb0gZGtfbHeVk0OEV6uWjEv0Q
r4jBKrMn58QuL4lsqXW4YWvCNpn8Gc5CZ8yVxZiZioQCavIWOoqVH3fgSsUzPUUycL86p1oNdYgh
vUB+x1YaZwodfxhFjRFkYeK8EO4lRUUIi1mJvVy80ElHLaRXbM1lzZnw3TKU9s67pOHUVZ9oPwGT
VM32XkP0QcfyLVKfylwdRiVkFlDSwqQzASytjxzVHEYhT7YKafxO1ULMBS8LbeYcPEQahSpjHnTi
SunO2mYEkBDni1oL1xNYNB7zvfOCsZIxmA3bUxw36bekkbMKgRe83Wtct5+jiHUEKrH6NBKbKLU5
49iDDT/hFwwApmBCkeo9rXe+Vn1qVphaDxyYojmJgU0ZbiMWzwrOEXfLk5G5j0uuJMI2erYpLN6U
OJ9fITScN4w56ikFPIsHO18T7QYDX//ZmOoQYqSLytaesGlS/4O7C8l1f6USR4kELUw58A9Q/y2o
oSKE5X5wazEec4VhtQ7CQ0NuToG5UMPk/F6tt8uNu7kPbsGDo+Efaz1jJfFqQ98PD/4HnDcNEiCx
tVndUkqYvCD3HfVQXZ5KxTV/+OvK4QHpOEBVnS0xlkiCt7iZjHCfO9iJ9PyGhYiTW8AV7fAgCLH+
tN7W1YovSgMFwbLQkxgDUZra12nLQFn4OlUQ9FNzzTr6R4vHJdPoKNVzAodEeRTc1cCniIccA6gB
9R2PzHOXRo1BZdA7M+csSEd2PG4c6HpsTB8XCh86I620a2Bd28mH0OBPOV1CO6vzg2uzTfmyGRCh
RMKRG8yFVujnCFrdKrvl6B+dwCzDAFQrbX1zJGgQinVgCmL7yjQlXPryk9u20IiyWCvqprGroDId
5rSJ+6XUsETbdW9IBtB+OOAx/NcyJTOPEenMuQdgw3vbouFpjeGyDVZrS2+F2WuRlBCbCnZSIoLO
S7hrFxWsO9KMK8i1HOMKJYi1EQOydbgrKMmWPFtlcNfZ2u3O0c4hd6HbDWFcas3Gyu4EhiydbG11
IYcD25uGmYSVgphlEwKKDf+hQuvKGYPqw0uU2oswCGMxutYDpZkWEGQ/RCg8bgbtmfoSbeSNdumK
Tsr/nJG3pVFzkb0IvXRB68wCBKkexl+URJ8kB01/iUh+QtEbcsPV9ow1QldcYhIkXljOVZgvEFC+
Ifgq+CRkNmmsLj+V1DzCnBTDTuigtOLgbvkBBMcihijfUQEk6JN7a5zhFxj/mrMeeIYx2heoV7nt
u+dMmX/ZCFrUrWs45SCkQ69ylPgYgGmS3Tgu2Nkyz5sjEv2kdJlQ3+Xu6ofxkYrp3dUbNTztfHol
IT+Darj39jtgZoMCUhpmxZ2nHpWLsZaZEMWLKpYHx2MO1VDXJ39sgLf/ceDjY4tNV0/HUu15WDhw
cV6cziyhe/bK8SZMG7gMW/QOzj4aVUyiut9qRvn1I7FU1d/hH84+oZWLbvrNR8fXScD8GoP3Gyz9
QwCQwqvalpWfF6i+7k1qQHhURMOdGjzbv3RnzCpYnZkFKiI3jyhtBn1emF7wMYy0UOSYQ5ZNkffv
BA7gs674N4Mrr05KKP1E6jBGH48Bt2KMqPAHckA2nryikHQhtGth9tz2gANKO7KIxTuDYiLWwwRk
TQxhNzTBV3Eoi4nEGbbRQM6b3OD95uw5pUKKL7VzN3HUoFl6ys29kYWjhWet2CNz7dHggQ226ds8
aaJZ6gGRDAetjkuI/cJLOSdSWzytk57ilMIJhPJtBia4gKbaWNKJrQC5V3OZ2eHVtEn7zSHsbedV
0zPx6g4xSANf0Ai4mJMu6K1t5+330tG2WvU/eEWZ9VvdLGeyv04L/h71CmwA2JoyvnddMLtl2FLS
OdOFSK0dGwddHCcqFxJOXi81TU9eqPruzdkBFgn891tbLNKUM+Rw5cel8HATUAePBMQqVYl0y2gD
nzgz9T0Rv8SF8vGgM0dvwfBPrYKiWKCDJZE6yGn5uYXZN+8649C2kZ1oyWIk9AIUUhfei1KLY88I
Uzwdp2iBve/m7AlpR1T4w2sGnuoragsAvy4EW24LbJE/BYZNQp2+ATOphdtYA6bfg7qjvwVYtmy2
sidSWkJKf31Bf1wGQxOnq57q/o5PfUTlB5TsRGqC8dlB8SoTrosrDPl1Gi0cWUVG+cXysydimu/v
CrWf2xO9GzDz4d+dx3VDQW/WYVHNB2v319fSI5bZZwPXb5ccPAqib6FaiEzQU9EnRHiRgStBzMvU
HEK/XPxhiicAbnqbZWDpyePsKsG3fdC7WV1jUJpZhkIo7VxSyP/6Czv+2u6zeI6Ls0NQ9AJ4IESe
vmIhn0VZlX5rcsCjGWgz4V+0jaxBtoGgrJzsomATYx5WKhaVk03eZMwLOThx/cpizNJq8M06ohyB
pJNXsP286AwEh7XNggfHQK9uRd3kxlLEi9zCzFMSBA5nKBDMJBKqd9mZ7x3XfptZ0IQROCfpx4n2
gn8Gv3P9iX02ZLa5A8Hr+cFBDypAXo6sWqu4/oM8QiWtvq2ZP4yPbo6kQf9fULdL2vAe7oGr529z
9MfJ5jY4raXptsSszcGPAwp8J9O/G+h64QHV9w/R7kqOMVc+suFKdILIVyjx/iWCQzYeNeP6ocR9
8GxIojfQWG2kbhOqZvHrkNTQLCV41/qrWpVaakfeVhEJZTXSm5AXNKswlUexZxxQqxUfVEljwpmJ
HA6u1lX+mbcAtc7l6br7I6PPn+hj6Mb75UqeXud4nuz3+PKvik4G6B5+8B7l8FDxiRO30nxxKJwt
nLGtGqlM0nhBmcmuZZ6MEFxx2iF4kaQWrceATm9QB8FlTWHzb4ct9p00Jwv1pd2Rgwo5b9fPcp5g
IWYa/6fdjQvdRqLbgw61JEK1H26fsA1RxiRABeHYqQKAAextnzpaUY3xsHghk2RD4aatS4r9GW96
o+hHAh2QcISAv5AR+QXajWz9mYm7IULSLYSlvYRoiMB9HzwjJS6AV0p+Mke3t4DIi1cNmhgIZwfE
GqAbRBMB5DMjd8CsyjzgrootavvlNZlcyAwDeQV8uPvtg+8E/YG6GP4kgocCWGbx+B9wV1QVocUS
aLWZZqu8e6E2KoilG1e/sFPpNkxvlPmEHXon4fzMemSU/pbCYNf4GeXlBKyfT9pbwHsHk+iIPrGw
J/YxuDNSe6Dg9129IIfVm8GaVuhQuYIJlGQBOmV+J802KQl62yV01N/DZAqgKvoqaB4cyyjHbe5M
X7i6J6ev2124EkGI4P1S6r66SM6bnJyHD7pPJCATXkBXnAQOZph4poWDOXVHA/R/4G91UkNNrTYK
7zuZh2vEB7TWxO2tC+thzBXixgke8wdkRvngFeiZuGbohfLvEG7WI1qGsfP0zm+fk1pSbqhxXPDL
Moq7EPPd810FVZ2Sz0u1vCJl6c4tOqZuEljwDQDiLL7a6/lOmfKnlZEQ8Rsx9LXIg0gYL9N+6mRX
bBnCPnypnSiDjqhfHhBXh+EvBGevuWiPIWCwecxumfwnpTykixS6i/ZlDsURQh+76C7ChlfVdIYp
3zFie0CZCSojtixoI29kbrL20no23Gm6gE75F939uhXGqbAQdV77zw/oKPpqME+UoVol8YTcWApm
N7hfsaJY190WwnNW5P3ifX/Sa9nnrPRgt90J0kT3Nn/tEPpbP2YYvxJEpYUILeAfxTS+oMK7Ni5M
nM3Zaw2lDI8lgyyrxmH36PKOaXBfAXhca46Js2Zk8P04dLrEJ0YVHfwg5b7sFffLqZqiZC2mEiPy
gwgRmP8mo0XE5593Tn66ZBi0VddU8cIIa7nkioYOZvovqj2j9qUjaE8KVnUef5hqHmpwMBbqwy7w
qMl243SG4Sf0H7wV9vKWg1fzuu2d6sBCCvobh+M8TNQuhwkV9p5NMbq4K0yPFcJwgWjDp1bbKbmA
lMBeAqtWncK1aCVs1ayjSW/5dwSvyEr5nnUnb8APDQZhvZhxEJ/it+WdAhxDoKUNN4qoDoC7/ERk
gsnKZt9W2qYkZCz9arLjjPPNGA65JdMKcsU40GaG0qsyuEtXRqfinAKvuBn9YAEZNcNqiQ5t2SRq
6+kbDBbGoax54Ak4AN/SyDOhHRmmyD9lCv/qgEyQjphZ/3AfC2brS8oGW2IPh4ugd/O6hUGQ4/jr
AU/TvvvpMMZDIl3m70GTMoeY1XS5Ynvf2yOQT3g/0k44ZUzPI/VN+Dnm986Q5UvF6lxYiRTzGpHT
MWQbKOCAjscKSfW/wZB7NHRHyDv8jvBVvGFoevtZlsuB3FA5c1MlE9UFtRi0V2m7GcF1QhPeifGz
tPmyAHYJ5fO08tdP8caZeSUygkeqInpfsb3aPK+MHjIM77KZ10RXcG+mYOxg6RJ+MKZnIZ1WbkVX
AAvciknX3M6MZVfJQ1eJFxsl1zclDzP1wpW6ul4+xrAeQHjrwNV1gCwxv2gyJ4MtjWwN4U7v1lxh
3cUkB1CbwUDnDfCU8sljNd1/s3kC14n/LIr9vlGWvCXwfrXGayQUKP4jSUGGDZlE+NbBEqohbaE+
t2Aon3g1MtkfgBujULsYJzLnItXT2OzezUmw3xLlUmBAXIRedKY3o3AzfYBdXLr0OBVdzQiBaW/g
TJVfZa5DHw+HkS98ijtqHeg6AgBIXGRqq5hbA2pHs0b1efi4mkajdugCyAuvErZ4N85/bcz8Zfef
wEL7ECyzjjpxpJ8q3WwstgxB8rh7mATAkrNj102CUsswM6UeS+qfL3zS4dIZti4L5IisWaqB7i9G
quShTpCTKZbsDkqcxFqxBANdiCE54hfqaV3aEa+7qM1VaMKfv5F8VZ7TK7OjBAWZa32dHZwKNgi5
+qCI+IS+XjgjClZJ3IQhc/gwTkCuwWWGVJNtBx9YHhP36tcKS4qngQvrljXNNIS9gxBWsPcdIWJu
Oai3jkg2XeJOwcfAdJvLQFSmezxbkCCf0VnpVxVomSUMwEfsqbL/kLgdlZpp/GXiqIdXEjgJRUAs
7xCksrTXNb3NNmusn8mMwLkRTEsfpNDPd99dQLwjSZgPwAdKLFXnfRQim/yku8nxbaNGjMxGiXIg
0xbvuTdPzAiMDxJC1puAlKmfiPP+tyc5vb4mxsRZYmiTNB1xA6glYG1B6PQLrVXQzg2FSCsGQc2G
MU+Wbr4xnuKuw++64XgshNh6CbFeHcRiIF5M6N9romenNHL+MZCbaXkB0N8yjrWmvr4FMNa7oNt0
k1UirkCl+h7yrDbm+wOMVqZlFMoMRGofb9nQyDnnXNCcmAEdPFDtXduC4hBVj2INuutoKVKmZc+O
G5Frm2VJrMp+CdL0NNcvmI1q4Iggbg6lxPBnfsKmG4ZMI5YIRCTntFyT3UkqoVTZ/Ft7y4hScdex
KU3bwNwfwyPWd3o9Z4WHAaWWCaY8ScGDlJC8dW8AlH3lPJVp3FqO9toxfMdADUe2WOww2FbBUESJ
R886s5MWd13wtrf86eQh6co1C97uxkvxhztc0+p/CPpjvX9kqb3xBOwPhy20QkNHEv8YJ8mLm62S
tkY4tnch+oX52aPilDWIOeVj+HB4t+UN2pVDBq90gtiI772LQ6mo/LBkM2Fz4+Dvj07gyywJ2SS3
LPSqUDGsSbF589cDFtr2L7uCFk9GUc0VcETfu7W7NqOXA0Tu89IaC6JbfnZASmEw5wnrpqgC9NmO
wMLdrj5LMwDKMgD3j9Saq5Z3j2yIbC2aWt4QZiji1k+0bn/CUYoHV6QOrplqLR3vehQ62Q0kaOjM
LL3oCgY2UvzUzqGe+u4gFz0wBIS306wc7NVd5it4WssdIbYoYRIGKVUbwRzG/JxcmdtNzd0ZV8ul
K7xgBxBr4IzfDGP12CcoW9C/HypydcC52W+Q0P+BucB5lx1zIx/b8azUNSPpOQna+Up2ok7teeuD
7uanQPl9CJ8YCYfLG8+DxrnGTUZw5Xcmhrs/94B6YOdmfnSB5ybgPXwBOJd/adNfKOKxbd+V/ysU
xgkOhPXp1SSEuBMr9+d7AavNqTMM/JWhp0L0jhy74HH3QwdOQWAo5bDgzLgtYhvRPe3w6psqmW+m
8zU+F0Oe5S3bL20tirZZbBFyH4nIPB2TyT4qzpskOic6jAwfbZ1HU8QmhrAmus5eXJ2U6KYCg7vw
E2f7Me4mQ1qOcUZOJMjsOmLoGZpymrIROanDHCV4NCvnp10PgJdPBq8+Yp8s8ZVmbskdm87UlyKY
1BiQ4hqw5d7NeMNdY3se+V3Tgt9kU6b+6YYYreTlUXYBfct67ZCbKXU83JUX8nYhSlEWXd8FNWGE
rmQ8x62qA0h7kXMS86+ITHXuHQIrwtbPM7VEp2afme20ZydpLC2hpDDYENeEAcMrh+L1f+iJSo7h
X0r4FRFzaFDM6a11WLikXmmYYHA8RaquCvdJbeiVkm2kAxhViNEJDo2viXmQIk0PyvnioSGEb5We
w2jFqMCJm9rxO1f9LUlLX9SWSarNZj58JjibaWvIcJMDFTIvpOUfXZGxDFSj8Pk3HH0euhP3sFwp
7+dUbFnHVJQRKrhb16kunZHr4gDpBsSB6Qfz9Dumeu7/5cuhjYegaS4iLnF8OR0oStmH1sJZzA19
m6MvtPtlGZShmz+D5x1zGmxM/aVbgFkhG0aqNnmV6deAcyjtO3IwxRQOsH9YXfe/7AqnZuIM74ub
pNSsZJqqChP5W3/b38J6DOTgZCUWoTDqrDY0X3A6D58heLf6w7EBjltm2wlIqMWmAn0IZwBMY22w
2N/Y2SME6D4bCHyYON29shgloGCgfrbFyix4jWk5Fld1ldZh7cQ0pSh6EFe5nkaD45tjb00YbvLy
G6q6978Vu5yf/xMx+wZRyDSR7ZQJF5/yKg9O1fSrFlayOXivciWhYdbL/4fK1a1plDBSEUsZJ981
NuQxbe4qWlSH0qrtNsu4GrclwrLot4sCfrlqhY1L+P3f+JjHGDWMSsMqTXBNIyzNULhpt85lTKqX
3rkt1g1OAOXoqovuhnfxaKwl/mDB7oUvdnFdY5nbt+c5QfsaXSuSyPzIeiY13wCTI9ChggOqIxEL
p4GLGWC3+mejR7NU1wis7R2acltuM7PGDsT37Br0Z1AaKVTPPX7OFYjOgBD4s7dazqiTmattfVIH
HiLZ5gCkBbU0r4r2d3PtTn7Sb635S24IW5RIqYfGDY71vI+VpaKYbHa5KNhcmo2IGoF5O/x2Wi9z
ckknj5YrQ1gayQlCqc5u7Lp9jANjzd5G0st5w7RJ3t8Mrf35cbJFxqOlZflt11QT3VXP0ELXuok5
TxINmyS2W2q+j3ndihU8IBQBcQz1AbbDUL+78EnUSIQYhKrO5FPZP+kCU8/HYTurzVe1pXMniJMw
LLwFWxpG/e6BvXYmfyKi0alWtU1ikW2cUoWyaKkzg6gHi5da9iWDKJBGe/9uZNJ+hYans7za0oEJ
kBpK/X02IO7ueHvr2eYpFD3Hkn/FG4/oAV1clv7pY1fDUWU0q+PUuUVYDvo+McqyAkh2glrMpdGx
tVKHRQqtoo7myTqUZslA
`pragma protect end_protected
