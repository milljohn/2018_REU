// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0.1
// ALTERA_TIMESTAMP:Thu Jun  4 11:11:15 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AhmDW0D7uyuIMGnz24+2+bLEhSMgZvDF2saS6jxo1HKvmPaDOao6hDDKaPrr8dwC
Dy4Q/mWog16itAXweNamNbPNL+g7nBRZH49faiIZKS71HWKWMnVZHv1N0eBAawyl
ujQtsXMfernqkOp8ZqGojarJz0aPss4fzlONJddj0fM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
ijLig9p5xRJrbQVjUb8FA2UAzgJf0XMvThouAqWrV8YhVFTPuhL+R4mhODyRcNFP
8wxRKcaGueUBQhRtRO/okxzGSmGJDON2toSbJTJSsTI7SeSGjL8jeiIJvW4gE7vx
LmVSPIh74AOfDevack+ruowS41ZJB1eZJxkCT2PjFhV7JhCs3s3cAbfE8HdYTZnb
tf1kUBrNptu1d8fwVfqb9W0yUiYFOXnmjOlG7ZEx1T/3ljX7SDFhxdYjWT5KPML5
+7xWU2BKfxaYmlocKbiCfB0LMacltnSkrSTk6NwWoHScFGFe0ofCLXmdwZEto9qv
qLIgfbEWeIXQIH7e0J1ZeEajL6bFK5gxR4+SfORJJCm609bwADzUVFyXVKJlrOGs
3vwCMOUXV46kodOC8WtTKkr2cV+lzj6iEwFYNx0/o42wRt0XoKX9CxpaFGSsiOyk
P7bLpV7r6CAotu5Vp9n4LTEZzBNP9jd8UWEHMVEikFsWLIKfb8/6QSTM24KTHym/
Uty4KQYlPyff8ddCxhW7EcqLhiyZbxGlUQNLUuLOp02HpmDwKLzUyNaTV/P9fGvE
UMN6Y2uTEOr8+mLmCloOfz14tY8UpflaegKE/P03rb51oy2h0bNT3J+UoDjAGY7i
XDf1esMzCvK/9gtZSPs1pNKEde14p0PRIpJwVAksNKHjw7P2dCxyzCiICpDLU3sz
BDHaDxXcHxm1I4MOsko99eKcp903Mzbrj1KKcVnOIfcKeRVdKGXqjKU8GHScNAnB
6d8Fj/S19Jg46hGTRcktYDqPUpN0LBCAvpQeF7Xt7sI6rqoRBtDJXsBeYzLjubIr
Hr3WlOD8rpKrWVKTvcs6Pr4gM9tQOKBVgX5bxGQgc9pbHUr1S0bl5PJ34DHNvwoD
oa5XNpA7G5jnWXffEnfAyQ74+nQD/MCwAxNMlEzLKCXvIar55x2o15E+6q+MrCNM
em6bMrqfaHrFkCyMMLJibyuM/ESYbrSAtJFX1ZMWYvl9GAyEpNxIdNiotWCwU3D2
yzLmBm3r4HepT79zaXXfBl32Ddy7ac6cloMmwT0ddBxN10Am5bPptguEa/Gv1wAT
GW9aDHRg8JxzVkeOTOC6L4RXUMMCjW4q+pjQv4UM74V8l2Rhlcs9FKTC+L95XS7m
yf7/ipHJGX473wz4yprBUK9qjBV07PRuh7pLhl0mHQN8jwyAgkW27pRiCvw8/Xhr
I8UPBUf4iTP44oRXoxkxGGHFdUJoW7pQXQT/9dgXxe5JM3ZODncdkIWDUwwCoNcY
xz1OpuM7YPMZ+P0J5Utd3LN3OvnchOHf6MjPHGaz5xBq3khEdcNnVR3W9UpZI7mt
HxnokQ3m7a0QAkEesElAFj1YNPEPhebjUVFspTM+l+1eqqcmGhvM0FeM+nxSrJcz
v3rIzXNJ9BOS2fzMB+0nZSBm2cbcO7etWGch8Vx5anFNZgVjAx8KE20EBk3vkpGI
e/7Wv72XZ9eRuO8hT2P4nYylbnKk1HIIMhU4f9J4Ho/tIdalXCsUXArg8GXLURIq
iTMFbIoEGO4e8ZzzudUxAOzzo01zfV0f5/e6MLd3ZveqG08Ul51+fEF2Gcf7zDoG
6BsfvXop4nQUD9mCPZhUSa3JzUzYxKBPMeUmLpJc5ks3/C6b/BxH4fI2kKQw7RzN
WCe4VgTxclZqm2MlnqWsdC+HwL6SG5PHbxTV6768w8tXy6YvRfJ0u5dRgYV5Mcys
QpRpthkFhg/G8krZnO8wmx6yTNdSZU3Fzo+l/U27RcVYEJ26nLvHbu0uxyqiboHi
1v+5nGCK5A+mCkXSv9ch7rarH4dFT6VzlHrSnaTO7cQ0vfidI8i0ZQOmXQVdWXF6
BQw+7ZZt8wShWTuB8hccHSGq0cpSx/GdBgIwE15g1NNWqFqio4l1244KbzrpD9i+
Q7hjEBoEEB2fvB4TYkT7yfjgWmSiIKw874euO+593DvFJ5l7J0ORN+cSJJSAoea/
XDaD+lN4LpePELe3qXO6VJ2pk8TNqqIIzqb6R9NhcAehZEJPXPYgU4VMzlXuKT/w
OGwaFhDKTvX5LH3UNMdCEg9teGlRvFkljxlvItMcDESrekv+WJ5ueZofwmOyGBYo
6lh67OCI3rHmxKLphKIPEdq7SNcaIK71PWIUUQVqaNB2frq+ijP9Gy7I2byr/4Ae
6mMx3qxBydhgGXPk4HBfCQHGcnxOcaEHMVZGBws900PqV067JIr2Tf6o8BQ4fVoj
OmpVNYM5PKonKpqNgKdMsp73gXqWVN/psVpeaVyGBMpOGWaBs+cg+TbSBOEiVsmN
4JelGkY4s12rk7X02nfR59kx4LSVFopquAxwEvZFy1W2zmV4b+ki/3y9Acvhzzug
iqQ8rrHmz6NzmKF2kcj6Frp9dhpLBlADH57UZEIhEfHvtS6oW1Mg1Wodrr9Q3YFE
1bzQsHTsPq5hzbO8jJWhZyCzQej7F/ijQMqlgNBuHyXeoUNQlotu3e4vXaBi5PM3
/H2j1g9cBmEphO5OyXMUUme8AybuB6CKNuJ+jUG7k5G/D2JCo/lqFSdiS5fsQThJ
nEAodMM4kKfTomeSXGLu0BQhUdKgG+hPbNEMU/iyEkd6EIG1BKhw8Gf1rSR1k9E1
h0Jl0xahPGz6zTvV/ba/FMKumfhthDolCqWDwtQyHI5z1+K9HAorQnnNretXGlK7
Mrq+QK7HxEF63yQiO8VtWXVZBOKFiM1g3g8O55qByRCvngJ1M8WKwlSST4IXPv75
7S8O/3DohISlLicPi/w1+BBJf1v5SRexNXBTilgSrih4dVUFbxJPP7Ptm9XaWZUa
40kpOl1Rku/9KHXbDSmBR0/IcK69GRFq3dj4crAeebxd8RNmVrTM/JNtbh7jdy9t
a3cNw3VuvAwrKxuux5vOn8cww9U/suacKfiTzIiPLdO5G1NUA90FVYEeMIiSrkFc
790xQd7CXu3lfthxeQiQXatYmoyTZc1kXzWwdrF5uWb1oDVX0e9u9+eMriwGyh8P
7NauYm8zKi6Ou8dIY5LagJGzr30NVp2fbjSKtNo0Hjs0HEjKL3xMVwUzxVLgvoLo
2sHBY6G+fY8btI34hZSGpdQNprsg0LMculJFDSaSfXfU8l4KDPJ/yhaw7okiUUkg
FHwyzo+XeVR78cj/txJta9jnLv3in40iNPzUpUcGn2j8wFHedNJmZj5ixx6MGYxT
RoE+jQdugc5vAQetnEiT8MR18Oh1SwhDcd8IePeJ7+B3I4UAM13IaI+sorW1eyIO
71h0R220OVkjLHZ9Ycp8WMFZMbWTodjjq5s8vyLChDYeyyGiCxyIZ3R0PSJUgPS0
bWR5zNbGkNMswzTzmRWfxeYJ0PSmWfAG8UbhiDuv9BnKmoB+yfxSRPZAPNG7VPbZ
myhFErdT/P5tAgXkwBu89v1x+vOzt5JWJH/4hgUDFJ/26DlGb3UQt+k2er0DK7F9
KTXv45hJ4SnE9UUa75KLx8RM+WOC+kSTrI4ygLo6ofmc34jvpwA3soX5GyE19qJ6
nU9gc1aG1qh5rCXjuG6FFqN/EV26j5PKtQ33LGXWQaaHwezEd5lcN8n7+SInU2OC
/YhPc3wJoGYimDZTvuSFcHhwrPJ+JeZvZICR+I9Y+bfjXrCBV5gfHfzlqqX5Afyg
BZOtus4b3lS+k+oXkFY24b527Ud1j6h5w62+OpLuytlQqKVP5r6QFnMNzIIaC46O
efQPCub8COHOE6pZqpdZeXzLY7LDgfvEtTKgB99UkIN7iyObFwgGgQkYOTXaBSxL
AQyxjrpZEc/8X5Tt20Ftz/tVHef9IXAacNWI8yktw8ByvTvrsbhW4Kukk80rv5E8
KkoRNRYTsJvhZRJKvALk1no4ZlDP5S7BCNWgVigjRmyYAwRzVtafwsj4CHlGptUP
fACrrdynQmWV5uI7UTVuL+Y57vTNo+QQOOuY09jKeluh57sADViPPOaRdLdKE4Yw
15NHIAs8leBcn4DbqfVVmh1trqC4KaeCGgXxCm/pGlDSkHdypmfTaSZAM2qAj8EG
qmzQ5se2Hwcsv7wMKRD8y7wlXsxBbwEOBK4yEen4GrRQmgmqumKaQKPEZXTzSgeC
y1laMwVnGutCa08m0tUUTlJHF4M2paX0wukFgQZ9MIdjjpWlH5V8iYjIrZ7hnzRo
dsLWpFVuiQAnxjEDwPUIN04U4vuVrPcouv+LpVYl7H1yJrqMtyTpt7abdyBsI7/V
1e8BkiqN1t/fhzrPmHf3QfhxAimcSATmTBUMLXo7T3Bw5MfOGunJUrw6AyN03uuP
x4ySvbw6khcOTj7nV6w0ffgaOjCBF+YZ1a6COF80Ghs/KeZA+zEExAHbdkVKSWHY
82VTTCP37YVkzHdl14Y4i/WaUT540lMmOuqDcQEagGBs2eEi4txi2Gnedty2QuQS
2n9kLGGcBWkeLMmJfllp/l9MkAYXkOXafmYrb6kSyXV3XiiJeHke2/KOO0penmrq
OWWSwAd9cRRaXdS4c49Lxkf+AXLZkcCHZAj63ZFobneNPIHZwfs4F94S9sMJ7mGm
9oBXXeTwSigIhAasYy9lcKlr0HHq42c7lO/K5OGYpECAUIUpYA3CIyvuO7dVuzs+
O5/LzX8udENJA4cCav/nYrBHDaAbODg7O97uyEPMowpBwzVg3p2zLZy/LH7jdeKF
155TDAOXLYRaUcggWuE+ippQekz0WfJT8zF1dHDOZLz2CVkgMN//1/X8bMWOCVlo
76BBDUb+6GN5Dj4IGrurWN2uXbeDG/VRefGLbCCQGAX1h2o8EIVYsp4XN9jXu5SM
iqFswh9ALnCGeKtxPqH6cixNikISaL+a07VCUfgh69llX18DGAv1nrpqQqC8vlAn
VTZ5A+imi8A9QIe4Fgt2A+jjPh00raKw8G6xtOpe1x1p95rmK+II2tzrIOzb7dcO
64JcakHRvmHKRcIAfaVuODQXdrlufCoZBXHxlmjmdM8iqYRzwZg+m47cnHBS28O4
jZw8eIe5nNNPlRwQ1nQqTQTt8jaDnVFFJejW1SwxI943miglfCqo4FoBvhhvhtss
IcrGQecMAoJsTldx+lQo26DFc/vFKb9osNz6yvUrX6xS8fhpw/YG/utSzr6WIUmM
APn3Yjuxmvr0ryyMshpiqxI7bzieiZ/NPGUWwJvVw47xyrBS21npna6JF/juVbpS
WqGEOlnqjK2mMcVMhtk6+qyS80M25XXtnsyN5pK9osF9bmUlm2r/56nJHjDGeMrF
e3vWYUjZ/5EfsMMQ3MWskD0hRfSLWhZ6rbbcH9veUwd6K1drb7auiUWxz3WCMt17
T1rDmtxcnZN/ljjsk3lVn+RxYzPWtQltu5c9d36jc0ZaTqM5Fw+/Oum4GdGug9as
oE6L4LrLUnJNGNxNb9BiVhMT+zUB6brqbRIhxMhQsZqgWHoleSBmzeBtMD+p/Z54
zTWkvjixWcGzpgSxI3bCKMDx5yJuqtwddbWd90lQ++7lm6fSIKEIfWYoFUDZiyHQ
MTI+d952S93JeYoxvE8XK5LDvBAqo1SLvtQPWvauXOPlPn5jv+1al4E9NPwUAf8t
3TL36Fd93E4sMTQHyQ9u517oo63ouO1rAjgEkzn0Uw+grA8zbKlHMNhHSKAmbPM4
jSZh4uxOYSQwyBadV0ySJnCCGpo58SlXRaClt5xuWnDQlqjzK8HFGFx5EOvTuH6f
X5Ic5UWZqXxTWE2RrZ77MD72tWI6MDMIzR4JPb5Yz+HBaHbvnH0/3ognFGtbHp2S
HD73LdT7lwiACTC4JISw7coAvGEfb3/yokFXyHrn36l3dwqnFgihCTwWntfWCX/E
F3QgWpJbM1jS4JryVJitAYqaswLt/wXfVP7PoCmY+190BKRXGxvAYGowFPQjIgzx
dyS1hrb3dFfw8IPK/QsSo76Q/MEkKkjM4xY7wKe2j0SVhIy21diWWVBs3GotJUko
P7sQq2ZESpxvU3X5qoKKID6CtOffwTZQf7Tgyi+HFvqqeUG/iYj52DmnSOu8WTXx
4MrL9J50GSwoaXTPwTbvZmAdeu/wLIPd3t7PGYwVa//7hgvT5O+5yj7sG6KjK9jr
R01wx+LEpISh0Tp6RMdcVnwQTBtAemm0AT0rM6NtgDihOVBhqFnjOBQrOVObS+RX
oRPBsSlhSjKQx8VVZl8825HJb6/E/ebT3UE9nZCHn9/dPsNB0Fd0z/QulH2/bb8W
/FBgYHHF2FFNvhoCV3egCNR/vtx7dRlAMkaNycojYnZODeLF/Ktw/yaWQa3qIg6T
cWuY9gbL8oc/CKgkMrMuJy6KB/a25PiyNZDcC3PXqKf8HO9hoWTaj0jbgkkaybi8
eB0Z2FqSYhjGcZXXmM3agsFxzMSHqCM5WAy1wlkAqSZ7WvsL9HUMj4/9T7EzERDE
r51b0z/kPaCZpPoHcu7kLaL4ptki7lQvEfmjIMJ2Ja7fKVC/trYk1zUPRAgK1imS
2AolfG8mjUWEpEkF14P59wHjECp5LCqoGeQIExCBTTeDnnJVA7D8G+Oh1nKnRzIl
vpQJSRMEeDozIGwy4W0nAlxbla8kkFqyJWTmcgmRfHfaWxtYpxvnha0h12EU/Lrt
6LJ/Pp6PoOfXODtYAk9gqL0PPrSGOgHpsh5JESZzs1+447yhWnqVxgvARHbNSppe
Q5cLfUQdSYqBy94Ka/lD7/luc/gzY5mglVgu8+diNZ1xdBXNeJO6YH9C55Y6iY8u
SIboHTSNbDIT+c2dQoR67CUgKfHY91T4qUv/wIIzp2RtRBNX/lhThJc0DmSX14Bb
HhLOdE+xHoqznW07MVpwKk0MbyWPR6yTRwQI3LDmS/d9Nyo6i+ZiVZEWN8mKQu0X
aK8ER31UTgNIDpMHdLn+9HSTa5ES40QdoWYJsQyPpiXkYMDCP9zGq1yGtWAuymMF
27Lr4IRCp6h9LYD8BAF3C0+45cjLDmawDpfbzQiOjQeQ3B2Wj2BrwtEy+a099tcf
OrNxkQRvsmYoCqsoayNESTB7UH5GlcZUYmuY7FmLg8XXVEtTEqRPdUd32TLvBOZN
7Cd95mdRPR9agybAIN4N/GzcdZHtXfSi7QDpNIvUMr0A166xBueyBkF5du8ufCpu
5QNM+alYR9HGzgKuCSk4+h4N0Na2MA/LYMqjyKoaeUXyeQMF7meWXZzugtm0iwmi
CKlDQtF2dBF+7i8oHy5p/g8g9/xr5qQOBj3XYTmq6go4OdUSSpXee736vnMVCm8Z
Dget4Gfty+ntMQLEEdj9v9CAxA98Ug3KblC4n5m8DxMFOk3pF0MPJ0Tj2ANtt/fI
9DYJR/UYU59LFdPmcFDPVLzsl61Eq/z7h7NHQu6c1Y0zC1Q/nuA+jsu/QsD747x4
Cv1y7gGegmQUEGRd/ZgMu1nUvcd4p8yJfaNbyDA/6KnZeKU0oHW3gh6aqzcF6S9W
/bJdvWnoKHMu5rxJzydPi7cMwQ3C+17+DfSQ2dYZYVEUQP+qdoJghZENM5kbSKil
z9QdS29TE0WwrsEPtvpe9vIzK7b2ZXbXWzyKIsW9rUJ1s6D74MespqA9eUsMNemR
EVb/67oIFLZ0/74vr+/mLbqNt21VyCa9Ehs0IQh4FXyvqZHc/xObhmdBK/N+YVil
deCaxt5MRYZidOoKrEE6Y5FkxMhqRYJCRFb5G0Z3HsFP5V2aOU21oaDToMmPyQra
mUhBlW/JnCSr8dC0Ry8aAMqtOYJQoUev13OWZgU2aU9EIMdAdfPk7HTy9ZYaEND8
v6ZPuBLvDNrOmbjv2bpee+au7aCWggoDe60I/+DLGbd0XAhZlZoOl9eyhqDsI+cg
PGPtyXo3WycwuZtM9DjQfGpqe45ZYHXwSk2jlF3IeifyDX6jkiwYaAXxy780DAwl
s/L13GWQknbf8Oe3dT/UsGQ3geuSacsVx7H6H9HY8qtm7aUl0kzNOjawY8mG4BXQ
3KL1j3iIBpPs0d3A5dy0gCVDRZhrxmFhTwM80ivNkpxGb0SljkvhljgQmNdJNyLI
AykgbgI6MRdp22vT3zaEnRyVT6oJAQAX8KVFdyTe4+KkLvuKDNPw/2rPVNNOg+GO
Sn8iTaPvYQM2hugHXBAalvUXTrO3FTHsluL88bGVbWKVpq9IFxSPhWldmsED3HZD
Ig4OX1BrCA9r0Tw/5SBNYqNxCyCUxOfGqT4lEKKQtNiQvfBLXQiNaRUx9DKAB4aj
iNSr7/uaI6sbBqhGbenPHQIOaiQrdQUfNEtuYDNrdLD5Y92k93KQlkk+rRzINBxu
R6xJoKi3z93Cx3oheMS1tIXsSrMxOx0rVuwyTr/abysIYaBsS+2EskBLzf1F7SoG
Z75vlxKWSnLGx34kAl0pygMSaiELLGaK//nB43guVd1diGIiIv6pJq0+PhltxD4z
prfYq2nTOBTzN6pg6jiGnta0Ylqv8kXDAIP65KVHThI3BaLEzDcm74/knIg3R6Nx
NFl0ES24tnl9ahryMJbBQ3I3K0XLxeaYbpVyh/fz0r7hJ3m6UNh9pAzy1ICV5hXu
gY/y0jk0c3vsYQql3C0CnKHUYS3a9UoFtbSncWfuP4rqiK76EMV7Kcuc37KdR/2M
Tzhm3e8nnRMQtk0RCqokKukN7n5y43WtEIznGTFkDoAcgSYLKpnHC7QsRNBxDuNk
n66oIn+2euUtCl0zcrWfvzY8rzWidvxImFOaNs7SHHdbbPrLabr9jlmkLDeWE0sU
HRwZ8++PyWi/PY4nfPf16BZa+0bjNWGSrRO/VyNVwTICbBoqeW8qSpR3Jr2L4HW2
AV7Pl/2FaMhvrESBMTyRwYhC9/nyzv4wkkGK+Lu9as8C3oYuogYj319FN0uOuP7g
wOPXksGP6VNnH3qakCIU8e8sAn0Q7Wg+ThQ4F75LxvE9/uYoG5iuQZyM2ZJFSO2s
1BO0sRV5u6QVX1Lx66EiUGS26KsRgY2Po8Vr6pVOcSCOA1uH/lZ39oDAPaQ1pA79
mCAboQvuhCrJh4QCHIggxFtNvBLPhzj+jSgcNRiuMqhGg9kh5OOEHlDL0tzYC4fW
wNv7iGqF9cmcf1gYYuTO6hmf/Ig4KeQ7ewCFzF+l9E1Qt9aSkAPk/c1hP3pxj/2/
ww5B5WpA8zrtBy1m4OdieJlx5w7se8T9in0VyD9P/iKKrYS/ikuDOughvn/PncvQ
9pjvVJYk7c1q0sDJD5RI/sLbXR9L+PQIccRLPx0JG5JJSCKCT5E6dSEewtjkfA6W
+XLs/pULjDiEmTV2l0X4WX94RaySq28XevzjpuimbH/buPL8Azwu4twnNqZl0xYI
NSUftqmXfRUSXB5J68G2TbF+kBJ7+/HCBTxAozAOfSDu1myBBdXQyqXUndZUagok
zCP3//jZn/B2RMpCspQTAVLpUXNpMTWqNuWzGq+Ac++p/dPbpwlNcnsdeO+Jx4v7
sGWpo2iBGDhgEM2m8Cn9+HA2KCZfsUQqa0t8kOTsYw3FkMTe37cNCnOrDvMQDmTU
TzqCnJFaK93Geztog7YcS3VTWVEATEUIUwv1s+/ZXE9UGSOtSuaHwoTJQ4/Dxe0S
n837dZub4ANZ3LpUFAXRcU7qHtpBL3qld+R8tC3HTyQ8+ydeRpyYnNawa4QbVK/K
pr7VJmQqpjedTSZcNXdI2fF2ho898iu2F4gpniM/UBH4fhucZHOFJGujcVwOxfEO
sEJdooiNr3Sf+EWmTdWEtI+qleY8iF6vMZm3c98Vpup05Iaw1Lb/gL3ydcas6l/h
qEoabFvebPGJprLd3Cp0Ae14wDTcUS7AXRwUNfqvXiin+AWHWkrKHpEANeVfaS/d
O7X1jEhuEoEWuVE7oNYyNFoYRhXWf4qe/QSsagoJvdHQG0Vi9yZCch3GUjYd3XNl
TE1SqK/63SDzSGhq2K19XEzkygUrjmuJvIz453MSZefAccWiri0WtIV0dWHaEM8A
Os5wsgpwzhEwyuyUrI/IpP5g78nP20HrSWlE3vDzt8UGmESTfT/p4ve8yGaNktQ5
wND6Peu5etBnNNI8yNJtpOkE0DRnA0x8JJOHIvxQ5RMj+de7tYvzRZGk+wJq2XCV
z1DUaddfs57DNsQetP2JCkfnUnbjOc6eGfH7qvHiuSDUknipuwSo0z2KqnIGh/CN
iKga7A54swIb5j+G+GlzF1IXNniY0QpCgU/5TvEW/75n+/jgJFQ/JqwUHTdZlOIn
/vW/z+dt8/XyHfihEwXZ0AWYPoZtWG3vBpXBGnUHdoTGEjT+/S4ebTmaeCa/Ia15
ZbU+TZ5FuWaSVCZ5O4cPRS9SZz4P7X8Be335wG8GoQZj7U/x17rVg9LA/YrkAzu8
P32bOGhWBoY0Y6utbSwuaK1gQoQmhgLukaOx1S7ifBZdGK9UXFJ1tBI3pccwk5zB
m+D4vSjEaljABD0XqIkubPenSNDDqBPSD5vRNOeuEfyi6a253Axc9EgRHAoxAVoy
uZ72gwWZmvpr566DcKOtOZTNQK6cwDKykAAVoMvpVAmDzJlThiPih95Zfxc4DbyP
/3t0yLPc/W646ak/1kflq3vnFMlPDVfEimRrOCPUdPWmZf+BbDm8OiKWionkovSJ
M+Tajlvo4+TPjSObVc2UiG927AF8z4XQ3KjsNO0CV8QgbWK+HsqHqWSlD8WwBeYO
o819D8SmuDObDhwvFMPLpDn04/6FgKGPBKxeyMSH6ZKGczH7Wc4T6V5osfcssIIp
rZwKF9XYqzD/ZU0KRH+SbwCFkWsf58a63eEPhGJrc7GdykVLHc03zfCJd2x40p/W
G1JchsBtcDWZ9ufNJDykOdbBPIFEW0FxyQ7UPcw2taIF3xDPnccsNWFqeJnxuhUi
oo47qAHjf2KMc1n8p4Iv6POv9j+/CXrwA4IaG+X6Wqmij5bIKahmXKItHnnY+/Go
JWE4NAKfmrO7fLOmr8edS28x69PDuLPsS9qdlknL0AS6FVUhXL2leiwFmgT0Atgy
pBHIiOWNlv0ZK3CKDjFCNpXOAmg202hM85oUMsDQRwO4vBE5JPjeFMi+uencmkTk
QV7H2Ny/1jtlX+ICWMGWyYhw0q0qqmOXluAsmB7/4kLILvaeKmJHPaCWMiuvL0Hz
fL3oee9f0ZEHhvp/ScorSmvpH247pNNBc619Yedlk2k21zMyC6TFoTyOrYwKlgKj
CcbjiLjDD33SJXkEm3VAaGmgpKuuZe+HLgTJcsoZUDEfLtxpdgL96ZZSoMmECvjw
lYJ2kWvHjDZZ6Kpugc2RJ28pXThUzKgZ3jev0e/oJUJxe+QAyse0LdII2S0KnNlx
JoZ9cE9L7m0JvHnrTs5ZjyJ0c1uzgKEJkEcfhrR/AvfWlkyspxE7mE+VbNbBbakC
r+RsrwS7sSOt2udvg83hiXB0mYTIITcAZKExFqyyRR2LyBua03O0lyRXunvduQ3Y
WgKIs70xzqwoBzZeQOwFqiNiC3KF/p+4/m4PPFrgqwddbDFY7pHeoYJ8IH3vqwp+
arADSkB8jjum0h61Ixfjg0uI86hYigE82tSBKql0uar/e2Vxt7HecB3EU53k1ueq
NO18vdtg6LPOREbtc3DCnBh/TVN1OPvlZK5M7eP8bzppmL+1zPbR2oQtF/FGcL28
VSJq6NZjNEH1sMZDt5hxRInhH+geWyzObFtD3+/OxP+2ABWid5996EFNGtQ9UOJQ
0yiu7JuUdZcXcD+/PdNBc/rjrBeRUW3N/mEzWPUPeGHu9DrjLSygLdIwS2Cvg6lm
GBKRexctiBTwEK/K45r9O/7J3E9BEDpBYiOCs9LpxQ89y8Cl7fjiFRswWZnopVoA
JiAdgN1/gb3+lG1zcDOP+XBdjQ43NtMxmm3ZufPwxRIKC7FRqNaoloLnKo7aMqPz
Ur44qVKR4q4F4+BAyMWkvxQAPYS8RTBnOx1wabMO12bzfccq3oKhJt8i2iRW0QOY
eCTxMOPTdNEDu9Zd1ReAWqArUEBKUh4fRbQY9S+nIeEyH+X5D7i6APUyIgOHMTbv
EUwV9zuKpgzJZ2xMFDYT7k2LO7ZMK2PXRopDTRglG3a5YXeNuu1ud844TxvQkDHC
UMFkaDW2pdFiPQeM3Fep01D+n+nJ9T83+TxiEzSq8WZFgAOzVA5pvjhNP1gZUrC+
eqnKOg2fIoRNzouRpv+SKQlo3GdwgW6mReKYEcYsYm5hjTBKgwkEvx8w3J+wdvks
wKN6/YFdXG9VpbzN/s0pNbUSm11upVMlsE0sgOpcws9G6+gNCWqI/I7aDfpPzZBt
Gi3iBKvyemkQlZHrZfAoZTmlgsDRZrI1tQq3aur1z1PrI1aCW/Hi1ENBHYNiFKfZ
sn9W/dRPL/LHC9dv0W8BXPz6rhrdm3x2mQNvgrJZq6wMVZ35WotCks6kYgU8kOWf
WSSroG9b9a17j9vtCvFEH4qrIOZd2PV2nefZU9KEbu7g000c8aP6sIzXskCQxhb5
TSPO5MLQJ66gx54uhegS6GpIUzrzO3MMyA4+oYFl/n/lYMq0bJyLm7R7xo+6ut7t
Ty8xRmRcw45Nrx/fy+dOLuG91z9MBU4NgejNVWtFQ0juRZ4tqdhTLLrg5o0jg5VH
HD+o8+IC7JsIY4MpQFzp2Yeyp8clFxak2Z7NPgk2F97c0R2nR36849BBrLjJarLO
it583IkeGWHkPrEQA+ywg2peY3gHj972bRxL8l9Oxg54GwSpTwW3xXYPGOX9i2yY
cbN+sxQsUf3kQ8TUscbKA7yYIhcGuSVVT/jRIOtA+XRKnk2sZiWQTIpA5k58hhpm
fBOB2wJNR+6hZbo7TumW0SYh+D/j4UWFzAu4VD5+s/7BBozevqHwuxzBqAtgE0Js
cIzyo+fcZk+m0/obsuAQP+z3sUFMuR+AAG89h/Zyt5vaGA72zSY2X6T4GvmUp6U5
0/Jw+JjDLOfRYOFD544/yiD2a520zjD84QLCf68ubBscieNMiWUFIA+GBtmcnSYF
ACwyW1ppRj6ACCSTwCFbX7KCo0n6HBLMg9MrAhwkmfFgLgVc4TeaeF3sc2hfXfoP
dCCYEQltw//JVeD1jygvV9AbPbedFKm+slc0jQ/3Gf90DhQLKfnZfCFAgxYzxE+a
Vn2AvQS9bsMBe525FpFkyiV1ylOdgMeEjmmxOKhPOGrp/kdvScti8yy1uRt/kPOT
QhSY0buZt6Py4hHVNWwU+62/eIp+Ku7DPyYNS+xLyt+T64R0VovqzlchvpjLYGtx
k2IRujuaGi7QqZvlUHw8glSGDqeHGMkehOrsFaWxG7AKdCp+o01YK+T/OAhGJllq
lXV44lMmm6HpOT3ZbUsu2Z1UPGvfL/yKgnTwtKc5UJt2oU61DMhJfno/ib8z8Shi
Lv2iDQre+usi1G9l85pmrMY33iK3HBdcwbgD8AaDG5U+zs2A2MfFSUxGsFO4U/f3
ApDtj7T9x622k5kWgIdTWlVinaiL4jfo7KVxBa7HN8Bv4DJAeHG1QzfeMttp7diU
BbCkt8i/EwmoanQRT1v+rYkGqW3dqgw5arP3o8fNbFGsypOqkG4I7GfTOqX+2iOE
gZd3aGanrtIuMSpYPRBG3xLrmVnCNs7nB937BytTCrqb+p4M8iDzwq2Y4BPkVfDV
VjwLzPTs87MsPnDJRunaLw8CAykgWNnNVtDCBSCDyeBO0JwKotKJ8axKzSu06fsx
4+Djp74izdvIwLP85Q/3TXCIQPH9kNTO/jyrXbYQa3cVsSLL00oMg7vpEb1r/7Ml
mUihSSoNF5eSeKLv+E6S9W17vtEEJLACCyuO8NGAQp214/Dlix4DvTLD9QSy9x0N
kXTF1NgEGZJvngUgHA6GjwC22e5Xe+XOKg1rlENO7T6kJ+K0dax7xlfC7i86gQtQ
dzMfL0eXCJmeXtQtnlBsKzkk9HF8gcGTcimVFbpWcV5xBjZ7so+YWX6AHV9jj9tw
oOr1BghBKxuUKkGl2d8QssxRuOHRgNr7uD9n1q9rrqp7sflRXXIJg0irEMNZRth5
JAP/zC3iqN9sHqok7oKWwv+4F+224PvLYCpgnwplZyMG/7nnQM+OGIdZZ/vEZXe5
/am6craAXf6m3AEjuah1Liql+397j+trDgKpzPnlB7Fb85Fl76cAAsBoMskuw2X/
RDv00RriOTYWaEnqD5ZaTodGag6d4gqqdNX3wtRH17wziYCfIOPShkAdUUVbI1Mf
sa/skdZUYz+LAH1F4vE/Uvei35UbvYs/yr3wcCnoK8wM0ENEnhaJnvrH2Wy6qE10
KJVa79yH6hDFp+EWbdon6VupO1Vi+KEbLovi7j4kDjiwf0EH4bvmo2yld2vq/DIy
Qz4Ynmlmrm1Vdup3qKmlfXzLkly5x8zjUaF9nd8Ha5vRoRv6QEs7xrd/AUkFOKW2
BNCqcnaQRR+RggGdXhr8FBz0btOlQVU1req/X9XAjq9EQ3SzMIxEV7QcNS4e9MXn
9p6lxsg8h19Wr5Id+Pw4fH+EohyJnESER9Nfbar4AJIweR5rGNAbwQwSrEytykNO
0zleWmu0VLMbcXH8EDb3EDExfl6qk0bQD1+AuqxYaMRal3kPS27zndMPTV3s72TU
zd1VRLah/crhLuoxKujkmYMCjm5fhxtDuvGx5Z4TPctNNggq++PY68QYAy19cS01
mTvHtmPyL7JKddtPFov1yl7juiRavqfQjjxilstbNQ6IIJrvB0rMv96AT00ZxEjL
FZhgQzNiILvvCp2VLEHpDq4lniwchGBiYg762DaaweRBJmjXHmYoivVYy/1//6Rr
J0NrIvwAPUVG17Qz7Ok0d3sD/HPYuxZxQRK0G7rA0M5LuRaoj7D446X4BAgOAy60
9w+UaR8u+xx4VlNbgrQXtiq2gp//yB6WYHNZP+Q4CxYWGHIu8Fw70Ylvi58a3Xct
1qL/LWQ+wpvo/aWKak4V3Oo6pKILV2/goNK+3e6XcUyJ4uHXH6XvCH7VoM0T+1P6
Q1qDtIwK2e+cVmgZBjdh7P8gWfnobPlj2rWUj6qABQ76Gf/KoyxFOlWRGw/8mGCL
JdjGlbqy65DAdFeX1w52mDA+kc7zqUK5O3C2UbdZighk7HeG8aHKbaWZb4DpE4vL
RuWPrAdnYYkVTUZkvdEf2XkcC+GLGfhmuOw0vCPW00DAzz3P/14f5PCHFuuegXS9
qnMbuHvKNNGFM8f+2U612AmYXZTAangDTvqpGPLhTq53oJs2XtCV/mT3Nz/IEeAY
yEsG/yGtCsZ7GswLlylDGOdOLOgu2bJshj+guspKk/rjqSTCtrdZ4HRcVhBHqwgl
rsQP/ZH0AvkxbPcFtaGV7egv1MygZtq4MVEh7hYPM7VffU6hj3nIMFmh9DvZuTKo
l2d6+p/CtEq6ZIQfuDm+ec5oRSSHsy95INvLGhAKNjn9bIGULv7JKNuZ9MRzS+wU
UIRHmRQE0BCGwKY0Sy0ZvLU3S2oY208Pjqk0c9rOWnIDrQKEDiCaH1RC8sR3dNBM
9AlmnJuCll5XH3nQ8nXft7XdruipsvF6KsDKv+W0N2s2Xm7eadpdNbBM6qa0GG11
G2GC5vwmcwDAk91dkLhWrG434Dk1CTRvqifbRiLY+M3bJZrPM+WgB8RHPGkI14Fa
o2pKET78Hl2i+P+MNy25OEC6iQ9zTGMtjhlw/vYkvXMvCsUli8IC9XqyBfIcqev4
M9xdqwYd1LR1CjTrOcnwQdoOSw83VVSkXXw1xCqnh6wMxxS5bgIUuRCxdq8jiUjY
RW2OyTHH16i1qmG46MaPROQmyXxgZcthck43zmRoc5ywxsI++mPvo01UN6NjR2wG
fgPbhA7ADGYp9Fnd5WEjWxN91VRVQAfRKEjA9qbMTeWkKYyNcQWr9AZmJnmLze4V
tTmiO9MV3vYiiElyxSg4Bv3b+WjsKWyXy0fIQC0c/4opPnz91Tz7sbd/YCBlbC7E
5HtouYpN2bdhIk6VfGw1ZLpP16AkPFQNVD5IrpKTzRrNGlTf/yyvaQzIBTqXg+/Q
UU0nPIgx4AvJPq1VuIjmeV6NPdqaB0JaguEzV9aVa3c4zqzSbf5CkeIsp/tIw2f7
y63HTufvz/9LuVie8WCpiUzobvxUI7CsbzeWBSRvTE+qbPuxf+JpXIClbFaRzv8w
ihcSs8J3gwAu98/dvOGSOBioXtcTtAPR+Sc7JixJhbI9kXpzaJYwHt/91Zvk6tfA
R6Ky5OjTjDnhywRmvdJ4ehA0YKrouV6PkYNJpo5OPjVSS/eT5dLhhwRVoRUxyRXx
Ai8tsulJgbB76kQRXDSzJXwQIZtQL5m3EqFvbIou2a03nWAS/WCdrDhgu/RKe1fN
d/nCuHME/zLlV/YAv1plJ9qZLADmPpYYhCr9aqF5nmLW6HNQtM9o7cDfgrLGiW+K
aCe207ihyHz6sVZ6URQthort8qat3uuctgTEk9XTJf3aTQGMqbuClJ60HW4/+6sH
DVkJVDnw0Usbe1iL79Fo3Rmj5n1D4HV2AKMk9jjd/V4QJ0DXSFceYkNLvbDJPqNG
Xl11B6mlW9VZZckPUv+N+wui3f1ScaOTD2N+7m2BgEUDeEdahO7gGQgccqApDG8X
25rjR9VC+LnXm8Ma231DbP1gNOI9lvyxagLsvUSViwzabqsBlgvkw5omU35Pl6IK
6ZmLIzN71QZppYCXs02Lr0X8nb+RgwBaolQgJWbZGWPjEjV+/K4kOALnkZHlDmEV
PNBUChRFW0mWKfZuBlVy7gkltZOC4qB3YUfmznmE44mqTMAhR/sS7MBmQBLxTb3a
7YfKG891NqbK9ZLXkuUbDmCfRTUfRsUyoVSY3iK9a7RhcaXgSBPYRvk+Oel0jB9I
FfR/EDK9gdkB5dxmg+EywZ04lykQ5GoHN6a/9v9AeXznlBFjcz/TFCGwS2dhfcZM
FdVyUynZexmForVKNjjSqf1kiSC1kTlEoC4w63PZMC4oYH+MVJ8B5x/1OTWvA+Rs
IILRzyJ5+3h7SW88Bx/OE4LeTcSMnLHr78EIV4ntvsID6QcpFrErE+IroPTNQ3o7
ApaDXyiXKNTli+NgVih+jIERu5VY8amLWQS/RrVQWuDW9/l0fXQDJ621Gh8gyb1D
pQOIIkhtkKYUzeTYJnfP+pAitULm0aaeqiYhLhTh40/ne/qLiVN+/dIzroEKNgUX
wWPGkvWaLyMul4SDcI7fxA56xIGGKXL/ufZZXcckqF48DbwRVBsKP2q3xcveEGmS
vIXrAdmXDQLN8a+2kKmabKISWLhgSuyWMYELGMipkQd8UNIs5kgXougsto8xQjOU
LgzRWozfGsv/kegiBtmZvlxrU4SoCqBYTzLDmO2MsZBMaV+wJg1k6MbkdH93ZJHg
1wqlF99DwyHFaZizLr3Bam/iOhKJb8tnCuODBimtGVJ2TfDMh3f/bp9W2pM/Tq9j
0tDDIK9iNaER239corql6f3TeQxDeoYM+OPaLQS9szc0WjO31NRL/4/m7XK+/4Iz
2Cg+Ktzp/CPXcuThMnC+8U1BCtdxYpBXRqpeQqJn62e+ZLCoF6xmruaA5v09Gm1T
RrGWwdlWfoGS7GKtIvhlKFg+GH8ZmDlL5YdP+Q2HDzrYAdLR0s/5aeHiv7KpgvSZ
cNseSiTRFJDs9To5AEnH40cVgiYZb2krFS0scPQMv4ru/yjco4Gsxki8KcshKqvH
fZC+YAZcZmCVqcNV9vNlZhx+/Y8dNcbgP2BTy78iEfN1UTWjHWkunIXQBD40fpYI
NWlmMR94YdLhG5INnZm5PbxgDSBIgmxXMbPnSF8nFK4EyQgDtclls/ZW5tUdmvUM
NJk77Kr0q0OYXR+Bmo8AZHJDN4A3Q9f79JrVY7v7+VD0FE9JJIm1JQSNdfwI5NG5
Qegr5ferNf/QYRAWEhxb6TsWDRllLZXbNrW/rhq/UkorGR4FuaqPs+7iPtJA7u5e
avB4z+482mGQw3hGHHkIB9JSKkkvUZgjZ/EsFND8GMlZLNqwofpCW0RLABFlRlKq
X9iqWeFWB+fLukvH/SZNzEQH22GrATbGbGsLwFB1jjZXTGLXdidET2+wi4cdHL7m
79c8hGo3UVnoioTao9ToyOBbsyZIE3zdyXRD4hO4paRR9ZTpl68h1SKdSNoSpyu9
Aap295oqhJsc51QukVwLXjFtVKU8tOMMexD6RMyFz2k0lCaVyIIkcGgfawc+asQ+
GzLkrPwKUx6y/qpXl+0e8CI0N0PL9DJmu2sUhWGfAb4GS9cO3uj3it01vlgzJsEp
+3vmxAugTl7s14NmX2gOeqGKmze1HteihZXxWjINjLAQgYofJ67wu9T8n1hAX0CT
UxtDL8tNBKIsmx50cUolyj96FXH+cm/GVrYBQLSL86MvpqZmSjp1ef25SH7rtfW/
TaZIPUOxD55xjCJ2mWgNDHHF5hyHad5OcH7L4SglIB6SQgp048Ha8G4mmDbuLGq4
VPmbG2l8BPRhqjGOMe3QJhLqe0l5zCvL61f3TSUI7x8ponpIPzfvJOeew4MsHD3j
0/cM7fQG/taKiOlFrVDG5FxE0I2m7nU0JTdvK2YGPihKD2VlrL5uQqUh/EWiD5LZ
tHDF3LbY1IVCKsF+EQuZsr/fIYw9iDHtOdviCrT5lissnkQvcZExpriEBDGUuZGI
2hnccx8eSGLEz6AeR7DdLhsscip8wQayzoVW1xtYcuHLyXo7euT+3mguqRzToCyG
aXKy17yRzLzzzBFieMzfqd9rQL0CShJAl0RBRxnRIqMDlaQXj2DXjN0N2kuC9ieL
dj6ceKmzO3aiWfI7dTwmBYMTmRK0h4t2uVmXtqx0uJMtCy999iDNPLGaq+AXOkdn
VCbU3J7iKfeOA16K+MFx0ylL2QtIx29HLAx/2HW4zkEIKSozSTCj1UIteo92PAng
hYy8MiD+H1zeGOLK6TkNB6toirT/UhCANx5I08XVZlrJQ8U8o3W9A1a0I7ESk/al
H7zlc+AHQ+XIqiRTZ8HoTFFgKBhNoTq22OL70X/BVSYqq71hej6jWEwyoBleJwns
mmMiEEZGfEQUINcyxUKXMvsCh9H/EtuRnIo/Aw1ERrVf/+xOM2ckTEm5/FGOlzcK
54wWBQVVPyKKjZ79WXhpRYt70OybdLtjkq7bTkYnXcL0LHMm0wUb4n8Qu4h3+iP9
WDe+tDOqWt9Yg668wBD/o2GwXXnTjKlQm+62uqnIpFlaTOpSfEWaG7/Vr1RVc1PA
mo/Eh7to+85sBnoB93LsXCh/Ip8w9hx2VVsTtjY80SFYjh6XKPpDOtxnKCuAw9ff
sVbRbHNCDpEcshVS1on87WM5IgpkzuKCBd/ZXYcdzVMXGOuGdkTvPJV7bU7cNZkd
5mTYSdymbXZbmubbkIIKl5Rpp3/sTtuMemyipuHKC7XXnqqpdHObqinG8Hw7P8lE
Bk+3cJAAF60UU52EcY4GeaF+HdDlWivqXxyOb7CC+Hbc3mNadEViYhDDo3W0B9YC
bMN2qU6bjv9moiari1UQxlFDuVYgfjyUrUFnx/CwbshDhwDKonnnRVPQ9vX+09fj
WWmQYBJJmyT3pA7AP2Td3tCdXaEXuUVI78OJnmb3z/9IUjC7zE4L5ywjfTJtK+Li
3bPzey4BXq9jqss4+Vkzad+OBwykfRl7J1m8Di11TRw6gLtLDR1AGRL2AfSCa1TX
VYbN8HO1tbXPdguQk9VRG+7jP8k3EOwyIh9zLRmVgl2/+9siCgmkL+9iUS27mQH4
O/JPIhfDzgFOgpw+3X0UxjvwWLgeNvJXTNFt1J5HbjsKWU4FffnhZVid/1WMrzyi
67U3LKn3FHiO022tOCLSKT72iQjdx5rWBtGN42KzBjC2Dfyj5s9jfPG5YvHG1bnR
BJ/rl2UdwRSbDpt54gmGC+E+jM4AabI0L4a5lpCfgAmzDG2r4kF9wdrMe6lqA7aZ
IhOHpqj55AcouAitkaJ65MoSTIXxPs+8KSpEMP3+95riAYiRja/ZpH1SVjH7SUkc
cy/ptqB1yl4OKXeW3FKx8oSyCWQIt8w5msbtkLO//J24UQW4WOhKF7HCJK3l6G1M
uSA4f5DzgwXOWDKwjo/xeXCy79OTWl5Qj01L4F+ALtmRMdodG1wwjK+SxVq0YhoB
7Pf8rF27eXkmGRMRJy2ViktSqCogD2M1MyAAqVMKUFCQJp9EHKw8YBsmrNYGUWyG
wdyY1R3XhYNOlrMx0ljeb0U/pwzlbKD4PANuqr+5rffw/Mn58N/EChccN3sDvCEG
JGyMKsM79B4TXddV1bhjxH5s92a4wbiaYpEwOtSGRi+TNqV3Xbohk1I/j6YfMsse
dl6pydZvL9nSlBSiuislPDdLLDAR5oD9mu6jM1wXRZiwfu+AIRIt7Fukz+G1rxpM
H+w5xjVyeOxdWwdW9nnm/Vu0qKYMrT977LY39JCs08YzHB/gxlmyDBG7Xfw6jFLE
RQPyqqfXNNyH4bzkwjRYPwA/kvauL9S1k36ERMA+742dhlrSkcCuxqfGZ231xoo2
WVrJdsJySkK8+dWOVScCdAYjKvnmZ/ge/lC+OexhD9TV9dwCvTCir17IDJxGE45s
sBxjteGa3AEE2UQrEEQaldyOdkAcx+rHpegklddd6nrcfdBa9S++MOOkL1/BRbpO
iXJKF/+JmcRyyi3lF4SBMPLIu+8Fbgqadf+Wz5OjSlYFT/0uGygJx0XPbba4zpzQ
Zw1tlwwmjMS2UtKp7mxOxU/lUpUyiQBW9TO8zMy7a+lEZUzsq8H3eUNV7vMipqUJ
WX518lwUvzh8vkeg3iOrDpk0GA69eBkIc56FQyUDrVHCryy8Cfg5vNrIIg/y/xN3
7AOrCwTLkJFo6q5q+KFImEhFAudULl3wbYH+DQwoI/h2IoRVt5ppBI+U8bJj2Xuo
FocxjLp3bAiC0xlAM0AIbAKCtJsoLT0dD0nA3JM29+4U55l/wuRpT+atApP93VW6
gVPzIHrO14S5l7+Vay0LE3HDPeZxszqSZtI8kQYrxQzFWsmnuoNpHeeO2kZlSdZF
Je0M2wS+84ksZv5GzFMzoR3kcyJ3shlfk6UxRr1sDYd4Ky0WjRhFgqDTiB2zfeLl
ArH4aAvTW+v5hM9jJtXMH1a7JwlYemUBbFqMnieZEUyc83KD7Ad0UQIXA6ksR0dv
zKEflYXA/57VRoaTv4kWaUv95no4Rqlfck7JElxd4em5cRy0EjwuTcGFfQ4bhFUk
ZaDy/19mTw/OmunwOVCYrds4xY+g/dikiQmBYrDDz2+5OWDj9HP9rnBxnHzvTggP
esNFMPia9ObA4ANLYLGhdMG0bv54h/E/kYPcxYkSXuwUvAG+vCYRbeIe9XqC/Dvo
llu2L/IYEx3ju3jt9pM6D2pG5Av0SnLRtyaN2TL0atB7d9D2MP2vpJ48XMX4WmYv
B81XO6wXwfugY4uSlYdVnx/E1Xlr04GeFjtVcWFMxkTtjuYCmq+T0OZvRmXV9NaT
WHKUXCwfgws4YNg8BSGkZlYR1vaN5cguzZWTJlcSXIV57LoaANTex+rR+9euHr37
r5P3RMJud/IjML54YCDA9Wn1fR61jyFlkbHWlitEEw9zlZ+483CzbTEZsptWkPin
Jr+9wmw/nRP3ZqxMeUECbG5zRzow2ZKYUlzHSK6W2faVsmGExA5/UiK42F13BBbp
DNmaGM4gugUpq4t0eMBJxNKDw/OkWZgoLNmO109QOOK5mIcBCCc5EWXAMOhyvNDO
74DKFp7aiuvDlTxyxF2eBObbKnuCcrblQUP14G2k1SdzyNIYU3H5Uob3dbb6egg6
q0JFKVMirD6D/iI/jJennDhO1czcnDFcuALgj4KYNk+j+rSVCOAs0ZvsFDb1OpfB
7YnnI9fnCEC5lowl1BFHnJ+0VXXyzzjygvt/TwKe9y7adBkZ07XjKLNVNuNDRKa/
IU1LjtdhY0lPAWivLf9ZXF/2NKyyoaOsufomEzikr+qO317mcsXU+xqxAGcXbkam
DDoa2SuK/ISD9SA6rXFCilEDqoelx6zrXutVBAVANgp5NCYRFLeop7pNlE/Ihufn
NxnsMrT3L+1VQ+mZ1WOFcmxtBA71v8+gmBO8u6IE6FKA4oCavZNJGLSbTJrQG+r3
0inYaGD5Q6nZmTLlUhXCnGi80ACrdIEQXyjEWcohUbMP6Awj+EGkkXDqD05i//Ir
kpc/ABf+UbOOKr2FCeB9emGiFuMWk5Xt1W/yS4GNbTH+lWIDt+3AVdX+i59m800l
jvifkHu3m8vF7tyjOML5M4F1kF6N/zW4Sa3uuSalTbLN+VbIISN3rZ2gHSDjA0ht
zm9xVZhv+Gqb6TjX6kuPah/wldFXOIWSp3dFvZKZIZqai/XQgE/ABIvsGg/8JZLS
DpGQVfnRsnvZTTymVoUeni0UfkI2DmEIR2vFM882sPH6+b6y3rWdPi19ayMY5o0G
tto8RkPHkuv2EojcbrhOTIzP/eAGdDEwlIr0M+8KvqgSgRPDysXotXeTyDFxRPWF
exIobT4dJ5PaeEJLOdOfczSgOouqGAI5epi92WUeghFgV4nuGWDfDFkod2Shp8Nn
erLmtNWszuVXkcLNnMuoI6ICCoftd5B4DfHBcQYoJxu5vdbvi87+aJLZuQxjy3GD
sCrjG18tM4BW7vHYiSs8uYs+QweZcj2sfSP47+WuXNiJBmNUZ8DVcktwmmrrJwNE
aaq+aNBwg8hfp/Zo3QhYC3+8tXrGb9FjEy9hUscnaaVQayMsmWkwxOEvMNmYbmOy
WDXoRM9T33pLyp1kl5SbU5tHuAXd8CmUev7CPAT6A3pPpOLViffAegXPqnAB9lUz
IZ5BZwgPfk7cbq0CgQgMzoI/SGA0DAfCUltxLCkGulEjCL0DUVoWeUoBewQQRdBJ
9Y3IEf6hiQA6ZMY72lDT2JUM8cnyIgxiq5/wg8ZIPiwB062CT2RyikYvDH4TmdOA
WGVsLQo4kyQcGzvYiak9xx3i9ElKEOgO4kGYn3o0mAXQJoHIJ7awrFQfJ7wf5CQY
qVQOJ08hI1V3X8MGHDJsLgsqGmGNm4m3GhgaDRfvLiWwLX63lKFuXoWlPEb6EYc+
0z6Z3j6oeQ6KOA5UqZS6UC6PBoOli5ELK86AvRgN/NtKdIlJeHMaXtW4gk65Xjhm
EyPFDi4u9ZDRcVhhW/CsdRYsO0LMpWZ5Iqt3z5UHtIsnp0cspD8n3i9/CGmBUzPc
YeqfylnhEppJEru20sHBB90LSSecZ3NDeNS+uOzcc94e7LkTD96t9xEygY0f2HLJ
WdYDcVLi24AfQ6SkfHS8ZbA5yOVEzE7XjKq6+4PQ4nVSMnRIXH9R97CWtIk1RNLk
yIFiFULi1c2CZuiO8wnMVUGK2OQS9HTsXTM6KEgDQt0=
`pragma protect end_protected
