// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
BPWHewEKc/i/MthiNpmPNY8uTx2DCRTC/rWuUjErWgRcEFbTfBC5shLNG2/cFLpWHP+IFFS+Qg8m
ckv4S8LtybVYOOHUPg9mjAOC9aJFWJYejTijSJnoIQtcchqSy8G0GPt3FcslhATpx53Jfa72m97H
dxls5oMckLIkXhq3eoHGk/FLX0bsX0fecRlfRqkUcmRA9N7xlcKCx6rthSC6uYzvvruce0XpdySb
bA6y8zy6aKP96T4QIAL8DoY/0ypF/Laj9FPQEkayKb1aLSP0+VjvgydXN3wwB/adj17MZ8PoaOT0
7vSz8oGN1faPkwzQWc9QIfGn69TqZVQ3WnN5cA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
JChbav26zgj4f+A2PAA5sddNsJstt515Q7j59FHeILJ/obmv3tx1wwIpDzQ8LoiOK0EstQkclBn8
juBIBd+LxW10K0s40Drq/c7TevNFDWFyFm1PWMjQsBa3MXYQ43oHrlQkLeatidM//OmQHbhTlyUl
YydL+l04EirDwBmU2GhD7fFMXSQ0WXkvLdZkpJyvPm7KBFrsa6tUGA10/gxkj47Afc+IuD0FoprM
4G9UU6ZrHVNGKi4/uwwNIYEXdLYpAeDWyPhZJSiKnU/Fuo0btM8ijKU3GNBkxqVjbX+B1hJdNkkj
p6FEjawSTFG8atzrE1A0pP7kRQ2o0p0VYNTi2pwQqHAOv7RBsW/1qgn5aL/C1plD0ylgT+1+U5Xl
SpfQf+3MSWutxRlpkKQp1b5iJvKcVR1L/9G5jIKTvZ7WC32KmfcOREMNtnh0nuiLYC7eC7jCb9tl
98ZcdxVWiIQFyNutc6tmmgSmk/dwo8GyLgTVX0EuR79qNGSm3MB/BbLPFcT1WKRKeWzD7ZmQ8S6s
4kl5ce4IgNPDkaS1B4iA+odNVFuooFjLkm7UVul2xj8CJzM8VVssNWPf9WSz0bUI7RvwTO/TMF5r
K4FnAflQEYeg2YOTXwgPrCQXo1oWdR65iOHZFbmLQT4SlxTLH/65KJxgf1zFfM1rFI9JcnF0fXaT
pyX7EFgux4e0Y9K7vW2d9rW4dMIfFdnnwxlOBJZqM3IHh71ddXykvPStImCFCcpd2bVgCR4Bysvl
Fx297chAq105wJdfdJNg0/8APUrGrhjzNYRvyz0ennPya6pHY/7PMNfSVqHr8y2RpCTAHuCDS/X5
PIF0yGnjU3+uXyMICSt6dFK64ckGIdtS1VtQ6lG8ZKKGI2i45ak4KVx14LbQoNs/eO4Qfj4J36oN
67a1Vl3IsoqXchmsVg7nv0x3RAT6RqNwdtLyhddhdF5z0Fv/PDh6sggz2NJQc2j4UHw47e0UNaGk
Q8JjwNcLLB8iC1gCScYENunZVwSCAehRCN+OnC8j6WSyrXlgEcffqBT/qx907i9Z50p85DpCd6Re
PqnQ+Eiyl2Cgi2PUQkzSSlLSrxB8qRL9RTelqEPIfotPG/gAsMNG/BtJiSLQAKJ7/oINoXfJeHJQ
FEHdec8wMlgcnnb57SsFr6Er5SCBNl7kiC+POQt0Z3Rd8OINDptZpEDXW1BGuBVaE8ioupzxopZm
sImMup+AxoO+SRFZkb5ZeMs8SjTz/Q4G+zITmHehUlbKqr0LW5bjpTjwJsR4D2KS7ClfszXT8qfy
buvfaZQpbb8v7bi9v9KPMZu4TuOms9xhO42FCTjsjo4LUwIiPJEd8VCcUQ2fuFik9kE8DWiIqgzt
sbGVIPSxF72intRAlE8drea+Z1SKDXDoYML92o6oWUzb4IWJzAAPeAKueVr/kA/Y2WQDkjDpBujl
DWcZHvRYgrhjGOH0onngBSP8vO/NL3TBmlpQDYXTy9MXkFkBytva04gz7r7pLLOArFzPth+CV6Yh
/TcmqfuWD1vcGU9Uwk3NU4i1t75jnAcTJVQrYPRxCBh5oMqlCTh+rbALI7r9ySxYwtcFmP4CyxJB
i2OvTuAcA5sDwBIK5gE6Wdph9kDQqaBU/dvjXfd/a2PrJXi2QLHN0zpytX/tASe2tq0bqio8pdw9
Lm5VAKjNY9x1gzq3JAAjbTa3za9kWhGbrDPojmmwH0Ivd6KjEtp0ouXbMXt3xv9tb7OryLmoa9B0
r0yJQNa8NmC8gDmqgoN0erXtnnJJ5vL10Eji1R6LUrr7iixWojANmot+ewyAgZCP6Ox4qMfQJo2+
YVPNhb0hURSsYXx6K+1Ox/JyLmM/8dLAk5NMVSMYjqxFbIGx6cuc51aLpPliCBgqbd3AYBOc7Kde
K0pit0KX7NkCPQEPJ5i3XPNLcRfQunhgz8nh+VdmcDZTaKzi7oXWtMhTpwh0pcoXW9hT3pPX1ZiG
6tuKNKAZZu13xdfmvb4fmVq72n1mTXJ3nol7CVzaTUVOMnQL0SicF49s9W3RsLPamSHMjL6VRueQ
ZS7fJyskuZ+cqoOZEdWM0tC+9QUBprgmJF8hu5/XlNkbljb/rtUsfY6Qghir9YokRpnieDakuZ4m
OmxCXNjnUphkptzDMSWSf7T38NXGmURc2DpkGM2iUKtNP5Z3QtOOHW4SFN7Dr+zlsOIv1w97KUTX
/VyoUoFg2f9dY/ko0bUhUBGWmltCYvOXBwov2Bp5+AHjZTYIKGjNnwxleYamm9ddCntoFMyRc8na
UeV36IgdV8FT0nj+z4RRdESq8mh4nKz2vIXT6tSv0cSoQv4bvv2RVus7sdnNSUDT+p+PfuVjl6Y0
vX/hcR8HLL63ArxGYesWiKBE4p21Uoe+ofldKYBOW5lYChybCtNNwUTEzYbZUdExFWKu6GSOPNM1
qp9WuwqzWu0y8I1kcvNyanpE7j54S+i/4b+jw19v2oRAm3Jc8mCjDfViy7rl9qkeVXm2arGMMD23
3+sUKYofp//SLkLqw1294kKV0PKUQIWhD6fAO5r2DKKwGIQQ/PtepN8wQIFY49Tz4MZWma6wds+5
LKesf/qraiobMknlW73rtGYwsbP4qQoPOEo3uwWs01Lt/5w6qogenj7nWOvXmG+KuGIF6IvTMxEQ
YUaY2MPIrdosIi7p6pYDxojS8wRS+DqshnZ5pi7QwGglVsWfz3HwcRD4+a52UAl5Q8I15itkdObf
Rm/A4KW8ujFm/Rqihz0XuoknIjjOEO2N/oyseW9kO/BEiV1fbyuaj6OHSHG0ph9brBs1H79qQ3/I
7M1vwgGFWvcqve6C5Jwfj0L4GTVIIx2yLEV9oIn5bhDqTRI7SndFGXQyLiY9IbKmoleJ8lH9Gg9C
YPckcgGifaAlw5WCm+k4wK/ZLpumjHp/M3nCV7qc39gv322ARBQBb7Nz8hzmfQ+Gxyy0msaoy4Cy
Ct9TPGSnjbutZHVhcZfZAqaG44nvxdQGhgEhLJcZLTdDlUmwpuM+tdjoVccidO9EIRULxy+Bfirv
PYevTN9uDDfgpe0BvQpetLUZFMYmVHDOGKstJPd1dTVz16LuBozb4uSO6K8itSvx41D3Ayi2+Cxt
Dbl6q12HKJQEhEHKn56a+Sf88fbnGMcpVm90BasLjhf2xlvkG7/nNdc6vlGcNNmR0dGrJqWW0Z9z
WcfvOOZSz6YiQ25h2vAxYjrb6/xLRQbTk5dF619w5k3MvtrfO15q885BfFujYskS6jsrGUvxo2KU
M8gCogZpboayNHU1Ywn/yAAKBTo+NqyE6yUGYLajlUnuNCbSkdwImaCaslht41Uf3PnfoP1TJ5wV
TVP2UCCFOnJdC4LetsA1jQK02O1xcI+PbBrUlBwY210wpZWbckHETF9OhsbR4RILkaZyPsQDzNx2
/4ybEE5LuuwWfcabeKMrbS6QGr42/fO66GUaTIFsLRj5e/JYdhcEP5b43gT0ufVR7xr1uRveD9ws
/gyr1YyfAul9N2N0/hUWroIyZtQF6inHNkabOJH4tCI1VYjuq4JscFGT/i1cUBgWmAtfrowf10Cm
Ja2RHTrUo966WP5rHYOW/EqoQ5Xk2oKa1PZ5sWmkf+9cpNlRBI4OYr/5Mn7zGZ0D+mAnEnWx0lq9
g7M7REcxKS21XCEO6XV5x/V7V4L1Qyt/yMkPuGFngyXYi02v/ubaGhDmcSrzn2gP9Q6bX+qH0Bft
WplCfW2PxHOHYj8O4aH2Uaic3XrtU5lG54oIv9IQ6DoKTitNTcy82P3qNF61gVQI1CT/mhtM9JqB
n6dyzIBttJ8irK/PCJ2JHHKjOjFZux9PVjVKQawMOVFk6ooBun4dS+54+Ws0Zi7PqLr0c+blFATz
N5ugXJ7fO03yiKsT7b4921UukwSbUjo/EgjqrN6XoCZis6Br+PTzwqGZ29ivUaK5Z1RNVyQb3CoM
0fDYTLB02odp5sjS1kRJ4DZeqRZGtaaH6PMkXYWvDJL1Sy/UFMhV82yVe9r2Y7DIIuxPi0eBgMBS
CRHldfuH4uxNOZGzhDE8UtJn8B4fJRDm0yOzyrLtkz37etTeftb4NMd4KGJMtzUPZjOkFm9bXdGv
QRMJBhARK9U6yN7nw+SiSgGLenQXZm/BE12Quu+c9gecGRDvu3rBEjfCzdZTOz1lGKzG+S/WauSA
CgNUcZCIwVGzcSx/jEJcpzB2R4aF7MvpbiaraIr4VvCb0LUjJLa+NAT609nh2BNzKLXb1Hgy+5xp
Udc6hY8bQ9K5aUCyx83d/5O+LNdMgaSQpr4jcg8RigM+gLUjefh42tdGw5NP8XU8surZnMkeHzvO
C4d4j3kujRWp7XbkB6TA3sb0+2N+njuD1CLhJ2QGY7X3dcidsWt8EaJGxJtWwzCnGXBKP3ayInNX
htJOQ2zOBd8yysBK6fFxtDU9PcDb4vZlDBojTjxwykro4qMhvMWNlHPjGjaoFYD6mcKyqdg8uqh3
RiBQ6xwLOrNU4M1xdRWWUK7Jzl3qdw433KFkxLfRsLEB3Pv57FSmAWdzh8t7maJXsHlrBRCaTKF0
tt3HnITxD7KbZfnqlxaDFuPNSZrQfDJI8sK8jg4ktMtEEZRF+msPtputlxpdr/CYy+06ZHvYNJp5
UHwMiI1Dkw6fV/+agYw7fth0AANTzz8H8ZuHVzMRaxc5pTFmehWdL0yDQd2V2XYAu9NUTdHFsqBe
1O6yrIwz3KBPFj1D0nQjcGzi7n7d47sq6WZ1sBY5+q8TgZDU8otNtzklV70J7Q9T3rUlFm/1q9fJ
GHfLBjIe3UWP2d6KfKDLSKT6aTCvI/ecfTx69YuqZ9dqFVJJqaLrEXzRgJK56jlwv0G3ZCtKiui7
RUeAXCrqNNCCRc9he1hPyW2X0F2elbjqZ/txcxf37m/RTskbohHHztOUHR0gGogh6Bcd/NPafaCI
vva7WMohOZ9GcO+VPW+IWiLB3aXG/QuDxXLuBofWB5jMpC9yTpNkt6whUerEcM27dBUhjK7h25Db
VUGg4tTNCVUDPUUz9QvRIf+qnWFQ664asnxBTOB8vpRgiZU7nw+srFPZWoeYRAcV+QXntuU3lT53
ug9vRFvRtx4zQjgwfp/Rsq+xvbfjMfHavNQn/GjYmkC47jEzfvuxqRBt6oEQpm8IYvAqwwGjw3DZ
S5lzm7tbVs72HNymvXz0KaqBFYF52D7yuC3iw4q4WTszD1pfN6cmxTMyo07qOSUtUtM+6UeVZNQp
E1kT6eT7z5HcYZAusnOc7FMfsouDAMeLXjNA9lCVoWRJZrTrfj3LpQpdTicMLr72nWPRKImNIdeG
pHyELZNVeP2s5QMfekVol9vjEFO9axcein/a7ei2PrJ/TAuhIG27klwRBZtQQHXGFchsbur/1KC1
9My+T5aOaXVTRoTTYvdxB8DDd60aTjnrJG6dcCzb8GblL6xqBmrfAgKDyOPaMJ54siUfCwucNZ/O
NGf/Ugs+YpjXd0WSLqYXrJiVNsaWN8TgOtHkKCibt/7rg/Z+8Fke020aU1Z4HxhMZZTbZDgBAawg
BBuXS9GsOMyWpWKAOKlvfp1oH7j/pINNQYL9LZcgS3AGENIkYiQo6fZjHCsHYr3DbxKY/7/EBw3x
t0lnUU4F+jCSAbRQKVr0YwjWDEVa5RhAMBVs9p/cMTmuLNOb0iuz38TK433MWDeMNMl72dlx2fCj
IPQOwkS/Pd8j7kvsuf89IwEyKeNj9Kf44DzjY25HlIhUmJQ89tI1YHiWDr9UHmyaLfFDZgs+GG43
fI7AC6vzifpCcAJrDfMYKTeLwCYl1kskCJ8qleeazpvzpYaEK20s0lPfmsfFuFm2cQv0Q/yGkBpY
qutf5Z8smsf5yfo7WV+voLZAPezM7A+cMIA4mI9OLJwK+ReLeP5TS88r5b6q9tBKSYG03cjD6wFw
T3aqnyuWIYaQj61yWt7Emx/BV+dB3dtjcZZx1L0aZkLJTBHKEsm5BLTWdH+fOROA5P+yFTx0Uqm5
zT3Hd12XnJGKBbOrMtjbxVUI/B3+gkdVovqFy2OJMDKjbhJlhIFMHj7WkPx+5MM3/oFhcfF4bRQD
JA/X7D4Lnn6KcvJv69Yfm9wOTkCJdUkvNBoEkq3F3rkw5ZG3SnRKR/wje9Tz7Atsk2x7M0fpSBfN
Ge2aPQtMALJwPEgq9R0O4xYgddcqS8TxTvu5O5yzHxCNt/8aAXa+x+9/ZPmN7oAFaFy15S04xAIU
/lcpbuzVOzPN1fY2ZwGUz/scwbaqrhVu7bCAi38XfOH5dy8mJVQWQ6eg32UuP39+C4TEkr7l37Jd
Ko615DKrnOt6jkZ46R3WpvKX12W8RwFjMiiHDyDeP9DF+rPkE04rz6UjdRcYpvjW7wafos0k/ROi
YLZZa2VXMISyAs/RIG3NCIukQlkr6UvB7hgvngKXRDpVWsksmMCLoLk0HN/Ae3wxj1qV3zIkmBkK
EHSv6IKy+VtnfJhOYvAlvUHF6q+Hawoc3KiApPxOBQd7XwqH/onwO85mhddDXCZJ++diti80e4xf
VtpJzaSRW9rK3ZVaHrZrKxmHRm49Gezs6TNe55cejIuiaJG8V6+6u3BhGC9IRU4Hd0UDfqC/d1hE
aE9yAtdH/fY7ZX8csuBFQUJaS3h4EmnxYeAgbFjmEQ/lqeJNtN77hqkvheli9fC89KfxYOcgCv2S
nDNrgthCztu7futtqwrjh64cG2Ak2XdCew8Iolt7RfVoGnzz3ioRbnwa4EWvxbzIsPEDeEP6ULx/
Zssm39XtzfUO5jIN3A6weaix1vExMaNr0NKaowwBegoJRXmaHD4XAY8Eqn+7tL4Lotnf7jig5WNt
4XfIG84ii030e48KdGgbKNrKcuq33PWZB5snaC/YvRp57E5dgRa7RwuF4AOC7QH8jt9Wd2d1wHmY
KX740oUkPVeoqGpzJnH9lnHQbSfbp0yNhByyfQb6lb938ntPSID3RYJdhFwPcm5F34PBlAL3Q9Mt
rMQjhSJdMiG0pOhbljc58EJRjZsjHBG8PFnICzSsgmFMJcWwBv1iXshXUiEAG1hRkkP02UJ6d9e4
lbUKcbNWs6phZD1856IeUmUw0P+NApLBczWQyq8i5vOpJdO4DHsltN0IVzmMJ5kcnJi5X7aZdqNT
hSlvKf8tr99AdgWFm07IsRcCvTyQElx51pKf0UABbuKpehhHe0G6XpIgvWhUJhxrZ4m7twDSQmWD
n+fivM1/3/WyDCzVryaLrb4ocSM8dFC1sVeoTjRz3ph8szRUxhUh7Jj5P8MtR7J1yP0n9N+VqmI4
wnpIXe0SNnJLk4VnUtRaT9qCpWW9LzOg22VZJi2E8hDnEQPoXc4Ja+r9W+BitFzKeC7FPTgsqyeo
UwZ0AliO418EatwMTwZpaWZsEEFzdaFfcVArWl1q8jRDJNd5b5EHp9lyWkpkJBdDLPV4Be/BrFu7
V5xIMxKAvcr5iVP7qkBWqNLIoD8u8+t2TCrEVAXYbjVA7DZccOWoIIIThnHX1ukEozlzirnFLSbh
xTs0O6PUFLJBoWEW3gZXYlo7obIynZFG62WQQTfdk4IWt4ojPS5tq12lMPLd4ALMQKm/UCojLaW4
r+YDXKqOURmEsxQs713a4ttmgI0ORF/Lsu0Zx/06CqAJsPwse8ZSwmAteM5/spsiZhSrWHCTyVhz
CkvlPaJvLi6N72C5pfwZO782ygXpoLviafdIfaaWJR3gWY37BjO3kTqyd+pjUIjqVmpQIwkzKX25
Rurev+vY4Yes9ud47nfdxew52F4mGOpEDLxCbU9O3HpeTAYOqEZ4E/pmRJslv6i6ENroezGMf/Uf
s/P43w6QRzhnSVsCyYVaBpz4KYceUsePTBvETg2fpHzEfQiDBiw/GCRBErqYTX1JEqw0rujW5N3R
vwe7GP73/v3JOJ6HDAXRsbQtAe7AwzSMjsaInsGrTuDzEj4yib2HScttJb/fFiuZapa7BhAz0l58
qMJUQwwHa4xqoYd/dAcPcOeRWsxAQsH3F1LuFCTys4/RIJgqjec1sAcYkuvq9THSdXj9HF3n9Gz2
pVZyYDs9fh2ZK7Htnf8R4TAWK++BPPa4Pzp07od87BO0smmHkjHnf979KJoGkSmbn9k1U3Al7vnb
QuhQ1D/7+L2EXJw5kxnx5PBX1FNlCbZsJpTFcAiNwgoXXEDf4QnXmwZSaJxpp+XlXlxfH4ZlYAMr
q3wzva2sUPgMNTeu2KoxnxaTsQOVCvUR+BUWbc6fPc8Pf/lz0GeIlCpk3MmtnR6qOMKd9R38eCkG
z1kCVs1gb5ugLa1HqmRa2VtDEXaygHPoaiqeRLaPlW1bg8Rnnc1uw4ZsqfRT78ArCVkkkr7Uyf1M
a0rrVLjjGbjb+q/WTQvCCrH9fQQaRBjBdkNYtIkPh8+7MFykGwlBAuzzlr9F1x7NQQre8Wz0D1Ry
1fgKa4K18QkVue4iBg+afHxd8yQxcvw/aS10cVTQ/zM/gri22GsrE6XL8pY0R5lWayS66J7Uw64t
JGsuRW1yp4UrzQX9GI6TJF4Lyi0NhacbpEk/AI1lAYM2/SEe2NCPKxcSr2UYxFCbLof97Sxr//Jh
Rkb0zULqSq0iKp4VvFmFZfk7/jQ5C1k24y0sEVPf4y0Rxz/3E5CV2/k0ibtzekbWUZ73PiCnLDuW
ZFFe6PYuEDP6HVZJ7UJPWHRPCAdCt7HhqPyEXpU6XLH1kLOIrXu/dHhss1ZdlmhLfkom/lnGYtNr
U1JYNmEeYreOocV1kFlN1YgEhzgGOppZUdJD+019c78DDrPB4N0NgTb6yvK3hesfCHcQPGIWTRVj
PomMUOFwM/J/0BorhXZ+da3/us5r5ZH1xDbjQfG3wc71fteSoLov1DfWeX6Iya0T/34rxR4M33bp
ZvdYNXZf9xTWQK+EA0FdKgdFbUbUZn6EcBXxGakzqBrsxZhuHOjo2h0YV6NIegJ4jkQOjxEqa0b3
kpfvQ6BMlxWxp5bfTGyJMjw4LoIieGHdG4/uS8uruPwIAwrZxLgqGnfccvyEhrVOXAyCmBmlymdn
KQmNHzNIGFhOroIkw1s++mwLJHehVAS1DBFskCgjUePQq1J8p9kes7kbBZVO8KoQhGknl8HvoeZ0
TOX9PRK1habdXDONJVGES0kwpodNU7sz3xlkceClUDpe6FVJ6YLMzg96IRropvOtapqJm/+o+1+J
2zW2CAh9+Gem4vtswX/mPFZWBdb7F3k5mJ83TIU2huINkExMjfuUtMDP6aDJhFw64KVgNYmCUBQu
VSKAyUNZN9Y3iEG2WGBYXam9S7jgNjBPxniIWXoR+YYq4JwuJDL9X0CAHAVgMV+OxWWHYyVYtDee
BmHfceAmOojxrc8REo4qXYNuyT2GJDMX+KuNuEfxDo3F9iGrXMBP4CLvkCIbtBtR+7/18a2Bh28r
yHXtWr0HWAyU7ab/0rS9eKKMd2K0vgV1jhqqvGUrhX4eA0B/YXKfkTvKRpnhDCKZ/wm6uTNhO1DD
Yy6/MYiuantjL7i60f4GWOrsjFBUVvCZKBYIjIebQ9d2ikY4ktdpYqO9uVcroXtz0nLDAfEPSfol
q4SxKeT3pl5fOA4E+yBA3SeS3/Kv0KMIsJS5DU40vBUqMEcy/WY0hAg51YffoC+ZzaZmGIwQGClV
4DlyO8ppVnuBt7osG9GsZA7oPsW9/ZtmSVQ6yMTgTisyJ4susSZ+P1k06IfNsbMUicmPFCXNkKzf
oAh90C28PO/2eiU9rSMNVEHmtYf8EQGaizNW5XZZXdIsu3wtQsHnxqtXu5Tw9yL55gKb6Htjtdhz
VeUx97dkyUPAv/O1wNDGxaIA6rQ/QAsElkqWNb3wKqngBeY0yIcFqM3gtaSqVNDH0BALhqQqdHWs
Od5am7ApYi3TloRCpqCus7oeJNhN3PzWsAK3O+8QxExTqW9Gxuf6eyR/rgWo2+iJ4kOZmK2Gl6xI
FrRqg0QyzqnB1hMnNukvM7Ivkxk/QSZ8Zmen6fjycPNipFftyH5jcIqdbz1ertCkD6yiazRcELt3
fwPtDLi0rNcRYTy6xdt8zkmHT0dT/CRCyfDMhFiWcJT1V6CbQxvCOwtaIHU+hp0iXFf2IpvaQ/au
wHfeo/8jWYHzyLfFGyEMky6pY32lu/xTyFQ8lsFzFXdsQJQ9ieFsW2Dch7t4zy8dXi7h9fO5kPVo
g7joa2hTCC2bqMQLveHCf4SmWBlYzAkZtYh+6GtNxgvmrP7OfnUNioIwBc5nrP+XeAPBISAu6U2E
2smsNTAJtevj7Z1WKOBBsRPk6ccJIt/nviD3d//usv5WyOrFdQPxza8mSCAL0R7hHtfOjrTw3+dO
ybAbtPAL4K/WVWvVulMzwY11XkKwapdA9k0hd1LKXfUrF9jEM1JGGevsDqo8L6JXB+LG4PKIxveD
vRF4ANtCo3QN3ErmYNnQKkzfwuiLd2iHI6lPvHjg9VTHfcDOhrZeMtXxaN0VSlLDAGhIY4S5Q9Lr
qVRErvPoIKghu1BfDuduRbWh4oqz8GXeBQrKzZ21KM0mE7S7daNZ98QARzCrWKfZEn4Vqox93Zs4
7YOWnpgDCCalOIjPDFind0aLY+rgrDi0vcLdar/9jvlZrGOmptARPLn+S7T+yaTlIg02FXGufOM3
TXxMGzlQtEZozBCLRjt0ebNb8i9KhskCviO63BcHm0UJruMFQo4ZdVx9a13doMlkBS219kQdHClU
NtwmV2yjwNzxO0ha3LA1YqzR9bdnvxyNzNK5UOeIGQhSqyZVB3Bt4EasoKKzeonJWpZ60/ES77It
8wChLGq6h8yS3dSzWTkkLhYKDUNEhwo7ezE9XmeHX7wL3I7fke/KxhVByoB0YIWzC6ts3rmviPAV
lkk2yICWQ05MwFcRJA1e0e/lWN65Mrn52hygIOfYk1b4agPFaBbFTZAnV9vPtByWGvP9ivAYfy1I
0YVE1mqPHAPxYAKFb8XMOyKS/A51Mjgf8SPPyiR0mjCLipjaB4t8pRkF5eexsG8cqYdN5gD5LpAA
QHH2H2AYeX1seEyDQE8xZ+wZkmJ3LfK/MTInVS8iP4XFW2hlUl0piHFdfuyblrfLaoqicI82tcvI
jF+8W029Qcg1gAPEC5gGuhUGEjtBAMs7dElo1EPegH4zJ2wRzZr8UIxNtJQJmFXhy+kkynqpfL2S
st+qUJvGcs0WvXlknQts4vkF4BWHHySm1oMlr8Yb6+tLNndekxd/HgZsum2LJcy9HsuiSIwa9PgJ
xGYuBwodFbFaQUgQF0llNk7b/8YuPeNCYFT/GUlbmnbc5hiIB49LXLA0mcAsWYReN63aS+xFtbo+
LaoCy2DhoQSwakYddOTNa4JX0MmF47NB6oqx2pG0cbonWIdc0IL+5kqHb5OAxfgQ6hIfNnjpk+mX
9ZiCAkY7VhEEIhx+lW02rJlGoqbbTSC0l3BsRZyfRPHB95V8pzbk/JuXLbVFOtdZfzSen7c36B2k
EsvXZsGDvSt8o6lrTtnyOezKoK47zAaDlgpLLVQ8GC8bmhnuGjQyWutFYPgyTFf3MQvQ0vt/7Sac
FG/CQki6SG+9Vf1QYu96TtaHKC77fOQKa3cacFd6XdByU5K/OKf3qu2pIksE8y5V9IXLffrmmoK1
BH1Oic1hZTRPBDquILog8rrUaFehkGxWbjuJUcEsVcv2m9ylQLcy0WIWmLQE5anrv/G8TMa34QSb
f9AcSXYyUSeZgQlBRJz1jmtfB0e0Wp5HZrERVtGkdZtV8K2gcvnKwTARVQwbRTyyRHuyTry8UcDD
aml6faXXeDQO21LBKFm/tXMFuFCTbj7YFAd3YQshWf3OXEOQsCFmoOjJaoou9p4t8u1CABPltcCi
F4OzqxH0z3j1XyrJkHpUgIQpIFGoH4B/z85nNYZdQOp1uv1H+ALDPSUF/j1K3oV7zewzGxFgfA65
OSo7OXHg+teSy3vUrHUdqwvrlwJ0ttt8sUPPMXbrakkFM2YD81Ir4a/22St2sUU/wQtO6TcCqrZj
tXhiFenJI5d4jJ8J3ftA/o7UbU0SuVptpCjG3McxVv33A3KIRLWeQ9QcASZr5nT6t2l9qJGtQJr6
xsQrIDocB5mxcXkOdrLnSp5zgjZmEZ8qclwQJpX+PKeWbedHnQRFikm/NWoYmD9wN0ucb5poFOaY
S2T8X4MCUe4VCTojqKU5bBWBkg9A/PjweXFK0sbqvcfnin9lFRt7RO55zfQNgAgJX9wBeODtxsLb
jpqPYC/+5NRm5Btpn3ZdORJjCskVa3hqPoZG7p1xI5ysqIsJAaoFDrmtu+GEazEjWi3ArdZC5xio
KQq4yPq3oNOZn6cGACnEZZykE+15O+EZPNTWIxmDEdCckXwaKv11fA2Vsepi6Y/GbLl6SwLSKRJR
hC3oMnojqo/62l8yiY2ccGtFTet7qQTDUSX3cwB7AQyccW9iUpvf2YAgIvEP8MnXjVEpGcVZlOHH
sBhc4ylbN6PfEERjYSLC6d0BM+P8Oa4DmEJr1aJDTq476RiqaSk7JBlbGUbDOw4P//ZQzVFpyOy2
TeCciV/ly8wKmdd/rAVVJ7RZ3US/9fT5QTB0qpFAXuV5coUfdSJM94OopIdQ35qjjUgOXTrPlvxp
Y7HBaWDFYmL77n+T3v3OLMfe3xAO9h4EPhIJeCAUVlFTBhcX6PT/D0e/GWHsqqDq7toBz1DYCTx1
1Hq0W4qRCJV8CGZlOcFrpXPgL5+BJpnHmC56UxtluFUae5LsP+HEi5inwX3DmpFJ7TMbTFwJ04i8
0T/CDXrJN/1/iDziApZpyYXGgo5Li9AovGNyf0qDSfEkO52PsUjr+QwH/O0X8A6z/kCRrqhtLYaZ
wvkuFBK1dFgl8eASu2D1fEQcMeDQOGrZZBDs3N8KmP1DbGSiqAfakEC+bicyDwmWB/pgswCHboOt
eKXfWtsKRDx3CDf+g7/ptssK1zIPimbROt+ZnX68BaaJdoUk2FfcIfkpTu/n3QN7jzPSvFqnlnk6
BguJ5cqTb4kvO/MJjGOfE5Llx4utVt4icnC4rddtBRQd72u+OoOHssng/7Q8hsXh//4708VWRpMQ
d3mvJogEif/JlEnF86f9hhXxvZXGQ8PZzdmuWrSaV20H1LKY+rdfDrbzsTKkZcIo8eSEEb5/YiPh
nhxDW6YgzmbJo3gQTSgIqqa6C0HCCQ6rZaFnronc2HRTWVmHGi6FDmZC3LNoMPqtd/JWeUy/ZeHw
Czap7MVLN4bvPXzohKUCVpZI+uoIJJtK5dthU34kZSV+zdk+g7DW30KGMzOblUYMK9a/jAV4HK8e
7vpvlmaQk0TxFgYptnRBhKGryVZcxJ5793kOxkxzd0EIEeiKGTlM0K9CjVfI1ExpcP4QdicHX7C7
IaKkHc375gkH1pOWegYCbnxXuiE24l1NsEoDMBNAFP3hiIUyWzMsYPTtLtEcFY2MH17HBEoXJnu7
BmtzjvjR8yjFQbzFP4+OEgBlCGe2UsyBeV9qhB9qrXpOszuxgOiXWhTHzATv6nUIJD22aucOBR9E
0zvv7BFIxWCUZ169j2Q6xD00Dl+m5Mv+HzAK2Dqe2+zv8fi0wfMvQpUmktXRKeB6KP2dYJ1YZMGI
k86whGo1Jtb6SmE9deaZr+5JuIpPaKwXHuwHTPyccR6+1XCeGmANDbQkuP7s8de3rIwvpM0+U2iZ
QQWBLVwMyq/JNsm0AuaveQ4BccUb1qse4UlSNrBhWmwObdYTwlIZ5q/3GvZJvndNe/cOGsfLY9Au
rvk8MbvLKIXwpGnzdYCOwQ3WWprySJ/e4INVz90og/y2ZBpbWCRrHS2yXN6kdMuplXH6umn4xc1p
ADzMd5cvVnD7QDGJ6xEtcTThJ3ZxdyJrL3jNOa2K3rDatugHnuOIWROQAyQ6xQY6kpjo9UiNonUF
DYmZqVUCZQck1eOHBdg3IdvaA7jZ8tfk+QHziB9hKJuv8bEAN9AFsJM6rQTOwLvZ7/OvS6O5kU6C
5o/LPeSTxjecPyEvKgaeZR16iCAxPpik6+senvS4lF8XyNVOWXt3Hnl4iRoryM8ck+ag+BaEPtf9
r1yX4DlGUt/PJlh0gDTJcJzA9mZchmlwMu8Yyt4ixnCAomJ0Pm9kXw5lKHlvlIEMTVvnwmN1mtVs
JIitOlXXwkgpL4CrpPPZ0X6U3PlJn8f0JVK2jx4ZZ1qTpzUIarGpkNG/C2P5JyHCLLTTGIgYQEdK
7BG9vg0wj3WQRkNgL5+UZScUrcDD8LjaYLqzTnDUbwtHwMXIDL+fz4VnhhKDwux5NVH3qNs/KDdN
v5Ksx3AGa473nPETt9UH8lngvuHbWag/YdtF3gagy0Qzhn3FdltBn2mVbSh6isfyxogsu90/URzU
4Ho31RL/xuA2sC4Ano0KnVJjasZuBn24gtv+prwj+M/+j1Fjoo/85ZKGeQ6eHCAvhTa8PdwME/f2
hAJHgh46hCl+eYbto8TmN8+xrr0yBTIZzWv794mANUXLX5yR/gaiAu5SFVE1rwWGmWxJlDo3Zcs2
g/hdjkUz8cwqdryB4fJjf3AHQgC6seOqANyBdWVNyobfQ0laknMJOtZxzZQju71IV/TkM9IAzOjl
kxzn0sQSCOagv6HsNFMwzLIuLPQpcc5WHqcOrjIiJiMDMcBIIU0m2BMm3+LeIwDBj3Lw7oCU0B7+
cfBYOYFM1nrod0GfFXn79ztr2gyh3KUvFuOlQARvN7kVKs8aD1HGDtyCg8BKoMxWy6PCYyIVr+WR
ahB7UVWzKig7DrsHKxNN8NXt42GrrCjoqS4TDa7r87QT5gLA5//xDkf+SquSGK88IDUEivJXdwdi
b+nD0PI90FCESf9bH9+EmauZTa13w3s0/OUvABHo15lA2OL5FEnQH0MTkTSiCZl54DmpjYL9Z3pe
SLrB6csmM9RTeddgiEp2YXZ8ko/3SPKjk8BcRX5kKKdDnybKqCWBKPSBUuO8dF+xEhTZ+xxohy2T
zus9bZ492TARmbHkafpe9Of+YlpjOuCFtbFHYUksP4DCbRYY6kYVyleZjpMoSLBz60Jnsu8Fr4NB
s+7X5pcshQBU47zYGbxFIfjuwZgitN6La64c49Th+wIE7Qhu+jxShX67scIzaXVrnW+/Un8dxH4P
KTnEV6F7LgwpA3k8qcNHHRF7vMka1p7KFPJeBKGPxbmu
`pragma protect end_protected
