// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0.1
// ALTERA_TIMESTAMP:Thu Jun  4 11:11:14 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IlUdEIPYDHiThYuIaoYmkPBldp3Lf9/hOfPHx7JcK8FqKhglIdBOa8ngatojU7xu
89FtBMbauWyE/P1sYBtB9dtWu7tOnH05Jk8OCErqSa0fDcJF8S+pj8v4BBVfzE5M
tVBr87bjd/hx97Mpq1ykuRXwbobxoN5VCZvvFsUIyjo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
MO7UGT6TnRCHicj/N0mWyOZm+VEAwVCaOIukQUsqk2hXetJyt+C0JM+J2n6lquFr
52jSnIvUP407+OaEzWKs18gnbBRI3xdaaCr7oinhHbLhJ2VBLFXSXwJM5Wl18+e+
otvLBy07rxsVSKMWUwxXr75sFMQM4FrdWI/z1YIYPl5HteHxmUEV+nQvSNix949Y
IoAT1SUKiVtZGA4wlCFjXcIeCDPqCeEYiWp+WhKsFP48y/hTWFa+Ef3pp/kRIkVb
9mL6Xg/uyyd5WvP8ErvOinr8HCpowS8fUxyM2wwlmZjn4F/AdhXf6wNiRPjzNHzt
fERuTREu7Ltc3tKr0eU2YP0tgDN7+hA6yyXoBHxfVOMIbU+b0De4rf21F9X2siiD
lzPX2BuZEe7wYm+kVAuE9uHMnYxAB/7IWMvCcmk6CNSZV31TgJCc8ZA6ntKU+ZFE
55PT+HPQJfvnaxnY0/i3BuRF0JTY+Xp01cv57bxLNh2OLSYBCdynNHndvPNAPE0P
PgaOT8bBSixYrOfe7Yqu0d+i4l+6yTrC31gR12IKkG6BISHec2yXGEVOSUW5ALPM
12pSBr2U7oml/WDM7hL4chLIJ+6s9Hpjeeq+AaANyyWuLwELFYq+aC/o3k9EgE74
jRwBAg+FNiCNeHcx5sGff3Ofo7bVeaRhE1DGWVIXfOp9t2sCU4SUA0ZjLbxcm5lJ
xePsxCGpvsaM58IIfoDoAHsd2bAKcpj7JE1BGzPwQCLqzzS5rNHbkyGIB/FWqbm5
dwuRU8QB56LEjFSrY9zfJgRuSFjOHQtyTyGDRgJFfpnkfJu8YFI9LupQmigjmEqq
HVd3dsEoij4z4trsBi2lySiyKwhuc29xPwSgctzRGDmBDF6mUP8fZPsnAe1SjVVn
UN3GJ4EQ7Yi5o8UGvgkk5VO3YjilyOHS37md/BRE2+B8Kr+x4JhjeabDBdQ9hhoI
TjsIJZauI1GPayJ0UFasOHefIOFJ8C7YnU4QN+9hOvjS3kvTzR5la4GDToLRGt0a
PwZqGqL7yyigaTHdy7CEsqULKi3yLv5mUFx68fErgKXeT29BtwWbDCJmXOZpJxri
uQphFdZ5QnwJPyo1Y6W0xpz3K2C9DkDkEmX7FEAWRbdYZllMJ7kOAp3qqPKvG48l
JzN3zcCulLrwoG85QNMMTzLpkU49RnFSnKBEYf7NVRIwgicYO661nqsf57bcrIKC
R0dNcBVhoIVVDvIKxyAMsR+Wb0tnpnw16gX79nzOJ9mxxxzVMVUAAQrZTdMpGkD2
Kdk5x3Vng4juETarThn0T/PzGQXBw6gvvN50XCCUKHgcrVaxYQwMA/jwdrf8EMuQ
ShzHNT4mdtrpJ9P77YQ+FFnBvo97/uyrkFb6FVsmt4w1b9fE1i6+1juWffg9SQ9f
uVAW2sqpMOBGcFy5O05hmfcs1SaJQcmN+9jPpKTYuV1HQs1ELFv0p/euBGyjZiRq
Qx/FYjTE2t5SfYuFwVmh86d1w1EyRDOZPngLX7mOA7v6gyvUA4nn6pkfoYbGuK14
2JRBZ7uTILuN760XAAzOJj94lUVlIXUsC6YGq7ENdyPkma6SU2zosHNPxNEBFyWG
LpMXlyBC2Le2uJCDYAhFaemWRs4Q9WTyTc0gQ3GHFsYz+5ScLEpfyA6iKmuqnov1
ckIGutb2BQT02uP5FBEWDdQ3J3/DmHVtSB9CCcszAMkGDNeTRJjMb73YwB5UnIf7
WwDIdinFtSfknIt0tKG/wLAylYYIlz7D9egWA9jfGPYLRqJoOjy9/x2w0EG0WMgF
k92UKqKnPrRSvka+n37ARn1RpHRWPyHPPxKr+6b67JFvUjX2vChe1u/SFdxbsaAW
qG6pYH7C4DZu1Ggttfxs7ZYHVrwh7olgOz4h5twSQEPTqNJw9Wv4PY2s1a8Q5Fvc
ApKHz59rjAArWSufRC6sAMbPxILAkQXynTcJjzxPRV1T28k+SK6nJGDqZ7/oS50Z
McoONc4HZfrwAoIVL+UR45dQXwdzh+LzXV6GPHpQlDAPE4kS2OeVqD5QqonrgX/E
uUPOn2iYccfMPML5h35FJOiXfXcQNYQ4iri+wrgbhFz8oHie0ZHdEk8+vQPFGi15
MKuTikREBPHndc2V9mIrT3rCPw/QnfEpn9DJCcEnxHSmfhgZE11ZyWFnZDGWo8/Y
Xlk94MmQvg4kq4JD918NMYsvUwnox4bGEsPz0qB69cwGVEff1M+T9sxEsMHcM2yO
Ov0ZRRR9q1us662Eq076YFq83YHF6sCqnrqg+gtpUEig/cN9AFPX59D8AbNUHCoW
KjZy6JGIQoRC548vFQB11XxiIDh6WBUM6XzDvmOH4pazS/+dxgu3vIVnNBmORCE4
qnOktmZIxV/NthUi5pacR4YKsrrl5LGbfHXqVSB2u/IfDzkCpxcNZ9V+rcw+dM4k
idO3fqo0XO2MPxgt7oVkTZDFetejK4SNQdYZ+HKtekrMBukljJtpMsDFCC4oybNu
15P44ELdnJc9qmX7flxmYyLGCeDlzLF5uLo1MIJ8RgOFjDoVFMv1liNgPRcGjvDl
AHEUIWeSgaD/1FuNhNo7PcqmHF1Tvq/6VZ/goYr89EAq1UJOJyfrpnHLGF+HBcx8
1iekBbzB2V8EHjs/MJEfNHw30TvkkPLC7obILyJB51gpsS9st380ZDjU2PzKMlDJ
uhfdKoayycaFIRj3TahxBbD9WKBpbou8vHR+GF8NrMjKpLR/4FJoRaYOVT4HrIiS
ZxpJAlkDwrTO711PLAtD7geeYLcWY4MahvPOBUGoj3veSMJUVzIT1K39/wHtV3pc
5BXs0INC9jlee10N2kJ0vxCZh3D/L67q5b8szhPCxG3yGQfl4ZAfMb+YRpwe17co
X8Q/COAhWMg6ECWpCWdURNyisErNSveLSkTUd7Og45WobG9+SxpImgeV07YbQJYg
QOrfkL02ANyG216UZKJaHDGU4+Blmu/Y4kJhigRCu/4A8ZEoF+dYdxFpTCadwFod
USpwBQ3t2wUWsPvcgZgHSLZ1B4yMs6LIlXzMDoxgPDYgtyHscB5x83FkY3nCk16U
ZvFnr6r9WE/KmJM13fEtfm+9L/8wv5zo81UNMfPSKADnfTNIpG2/qzCJdjlxc3jo
6+iuA7iwYNVUy9TiaY1Jr7XuttvGz8Wud35LxM62At+TGEYK03BGTS9XMfu3iUff
T8V95MPtiQiAk/ywmJuaHMG0OnIxn/O6BuH7dPZjdU5zus3Wj0ykLhMwKDLEOBWD
RZagW8+UdOjvJsMznW1FzxN/ODJVFlfSwSo03GOI8lWPf/O5fya3dwoc03j6qc2h
HWEK6KOvl/35wGYUVIMIWZLIIvRNc4+Xm5ew/sed9XC4OMGBB+TN42HZeCbTX0k7
oVYp3PPkmzpn76cKq+G8UovsUgnRw4PYsN72azeP+NuknXIQOTSd4U+OnEBj3lq8
22USwO6if664qeip2vdTT79HGlmHfAP3C7njvv6bJtIK95VUpWakVN3qhFnZVPyD
tvPlkTOoVjX3Gy81azRCNZBJ5lUYeQM1zA63+v1v4XHO82JKIoXyQzLe46kg+rr8
psdjM4BUr3piUdFQd2IG01vmB1VhvN6D4WoIdK63melKPGZWm/LOYRlp+RLU/dSh
fvZQJFozauWhlde/R7JKxsDQxisIPT3XWdBdrJSATr/PyRw/NdPIIZyTi81oWkSS
346JvH0WfM5woPG4J1ItxhufLTmmf2q0iv0R8AaKrt9ollQCPP/jmJUZfUBFmua2
8jnm9qe45gEnlnPjqRf4ct5coIYWkDbYvIot3sUESBA2CjqahfBI9f5yxrutAQgJ
e7Xk/LB3tF2IAo77OhnK5AhHhIZn7pk8moc6QbGzPiN0mc3WYgf0b1fOgrksBzAr
RR/0m3/deuYcuOUndwsItaEUk9Itkgwzo2GMU3rA4LpaGf2ylaAC7T0IEFXdZymb
aE4uTgdoctAPDBIoAyMZ5qB+BHO+8xxa3kYZl6BX41HCmucCR0NElLaW1F4WDLpb
dPP7R1Qg1o9EorOPZtIxEnWikGD00Tg0LZURxnuPQ08kjBmBJyx5XBsSMauEn5KK
UqIzuCfU09A6pB4Rvej7oX8dgebogT2D9j9k0gx57C8t4ra1Ox4bkCnqXGKShKwt
UCqYIsnL0ZCznDiZ7hsOIvoG1LBo97xVppRkngq+TO9cAD7SndJTXsPOEYKzdSvI
+9GgGKYIvXg6x//G4M/BvqQvhGTlj66Uv719f5dYClCCqgwiASb5D9QV8WALw3t4
OrLWJ1bdd7I0Nc1/wacqm2lXoHD6vNutc9BtuXmtOwUlqrupnUInzBzplebJ4e0l
gwPao5cFluy0Z6IMZk5Mz08YlwjNNpnEUQ51AQdVMUCPbWgckvkIj8Xl/uBeDGzL
NnaOxxKyy8mfAJiLSF7BJxtND8xDj+iRVZmiwPP/8V2q+5YXtcUWRmztYlw/wnjW
obIfHNaYGwGaAHDlN6GLjK0wVnVxelIa/Msdy26+mHFCKjO9GVm1O2fSNU8pNvUs
tok5CWRvAMftITzRKk8DSYiS6DLGHd0r/mOrFV7YaJd/BAT3N83tWRrbw/Qgp4Zz
0IL1BstLhL7LprDSTt5NssnrDSEMHLnSd/fBtoCNI07qkLIm5r9InJTt1W2ZPuzs
+cS93Kbzg0IatD5N0BFGRWQrXLjIBpaAXwIf8RJd9ClUx4PHcJsrWQqPZEOy0ZsY
2Lma09r2vg5woM9poFZJ5E1kW7J4zEi2B9CQN3tX6yFpgKNGA/CklupNkOsYPX5v
NPZShjsKMFP6RTGwFWXcMU2w7KLnb2MQ6xWmmFexhXvqv6h+m0AR89oXL4+Cl81X
KdsRYxajAVUQYFnRpwXz1x3nO3oub8EZAYMg+332LMNwcRoaOEwJ8vuvqLFCRM2I
Ykwnse3U6Z8JkedWMUMAQ2JgQB/HAdRoKQl/Z9w0BK0t4yzMseiPuzdOoAY8kYwg
hMlPGWUqoBAQ5/EvvWyjeCkel5MvZUj0xPoF05dzKh4dAwfTBph1ct5dG4r7HZ0N
WrNrTWfa6ocQjapyzujCZ3clBn1sLjxluc4xrEIgYZ84VdBE3wVgZ8CasZizaXlm
TF3zfKBd/HzKURRJAb57CP7i9z1xQ9V8l9kQBDu6OKzR0Y2Mi4FSlGm8HCeqj8vZ
1jD+kTsOX/ClDKyzuAB9jxi7rb1taYk984aDiweo0lXamIauS7ImklLHZAiuoVNI
PzUzXyIJv+JFVXUJlzRij1BoaOxr98rN1bCO+i1pVErZTSIbsl88yYSzr4Ys6aQQ
BKXEjonlfMrgjzFOfKQQe29xPR22sqiEN2skm23820yQSxCqN8x6TEca59RgYu7d
ws4KQhLlr+lYBVRrNRWYGl96sfaR2SYhIzo5/ZrHnhV/e+FOgn1lCdTlqtkS86OJ
NdbmKj3pm2w03FIIPjAbsHeeoih33hhqEZT4wKEoDM3pYXDzUobJjpLpl6eXlR8p
A8JdDjYYbW5pk0YqOtbrlluBL46A/lPpn6lDoHKE3Qo/ufdfXVA2MOyQ2oMhGwgr
E4d8oPZF/pPxLmeUohoC7lY1ygG55FqeFlptLys5HLZiGpuL46Vvzh1CSXsKFAy/
WM39YXgU5JKJL3MkkKckWko6xEviFp57DuvtiAaQB20A8XNs5hQXNusz6l3px8zp
kz5eQvfBZfKLaKcjA4Ey23mIg9rC1sIgkL5grel7j65iwQHGj+W2UHCrkheZmgd/
8xz/lk6lHTnL1G0DoRwfH/t7F33irBy7xP4TKD7BxXClfoNT7OkHj0mkzqVSwCUC
X4Jqtyg9Yb2aEt4h1oexqw7tGQYJPaH/77TMMXoaW8hVidTnSD43PTKHN0xyGEpo
RG+JyaxqPCYTyBtHgNUa6RVfc/0ChqanLxOwU5ByVRwOibAvzRKRaKbS+Ga4T1un
aiPegugHUGobmcb2n51i52nNnSQ2VNHFZJrmwoR1KDpXYQAva7EmUYAbG4WwMr8L
GtV3/tPVXS175oxpVk8mZz5ll4BkJwTz0Bw047ul/NX//DYIbYhIAwO63HDE6mEu
13cCe2Zwsq37edDzn29TSGE/DkiK2PZMB0w9ik/NZUv3WTdQmsqK6rRrhpbqndhN
TIsRJSiDWZPq0hAVhgExnkCzpGlxcKbgofU7kiTJJ2rjoVzf/G3RkDHfwcbB4nnZ
6xjFWG7vsKM6DXNZDz7Wc5c2jA+zsT326Sim56Ty1mo5ZmBayP2LSbkwV/Amf3hd
pYtUcBtf9D23hvpdd5Mkj3sMg1TDp9P6MZBLCDj+b5i/39CIzRSRSrrWXN7+ceXF
QKeYXWg/didd7JqwXHC9fsS0Fzk1g2yzJR3vRE6YtRfO3esgoTdG5/Wpy/pv+R9/
7FblEr+71WIeJS3YiCpmsWhg5XiAkUXwhR3Mnk1ICMIOzpTb4uUBJTMPKh+9h1Dk
5Olka9DBDe3Aybnb1DvIblHnyxvDYisZSWKUaFhje0HUnswnqeL5X0vEdht848GJ
CB5SfoXVCzhjikE9AMkv5bgZFpul3f03ijchBx/buqKSBuX6DWYfZpeK8Ml1fpo9
4Ia4XFE4x5eNrjHllp1ZkOQFiyR+IDYJg+X2nmJrB+xyw1ALoGc+xGmXSmTzSfZr
4f4GINPKgSAgwIUoo0m/BHMCxOsrRcavQGrNOWtlQMbQKiSQgaeddoFSgqwhTA9G
bQUrn0c15NeKbCRKWlr6B/s5UzbUl7dclEbu3Po91Hm2fKGU3Rcjn/Thntb93sLN
SAlkeIi9pHyMfWJgrTubTL1l360p00KFhOHsXsRndpY5PQ0dnT8+8Qc0YU71PDvp
X0xTNRw9k/YglSfU60MaWADOIQVwloPqjWFzy9oEcngpyHp8WnAM3HgLka69MYCS
y4sTTo+gQ177LbOrd8ELv0DSRjywNgE0GRY8hupGaTRHbwrPM9p3avna/fK8ghDX
BLKNH8etmzNJG1WRLXI8fcvOnYx54FpWdRM+x4y8QEuwPxmxcUO2cSwzvC2sEljc
ASYzh8LP9foDx5qzaxx11E9PiDjPtmf4I68GecIP4OPsgWxoKJerDbsYJYUSS5OV
xYUe5PXMHs1qxAZzYIrIpESgbIBJoPe8EdQSg/UB1uG1H/kYODX4TFqkRtIZgyVs
hD591tiWPW87UdpsCumeFCBQTIK+6su7swNC8RTT8sMsaTKGznILw5Wt9ULF7Wpz
GdJM4jPYArgeCNyDzvYEQmoz7I31fz1Iw4bHxgnE0U30v4DK7PrCjXDeee1LWvj/
ApwCSy/HHWNC+IqFFxTiGKS0NhoONWvkUaoV2L4QStUiFLJq/fYModNZKSLuZUVl
/UOxYEyenpjW7sQG+56rFxUd/Xdq7+DtnDrw1A4gbLKpkgq++zRLMTgRcHVuzgKy
+iVW80kb+SQek/1+dq9/SxChOXheTPnzNwMVOdwiAQQHNWBRIj/QIihAaknlD/y3
9oKCPiDzN/HT4Skj28/irlQmbO9E4ucarewFTQ2EmrugqXLkXAWFflZyry9Ebr1h
gnucK3Mq4w1SJSN3iet62I0SKxOuRcg71TwmFjVhuWB4B2B4JptY1TBwl3h3nagP
bJNRatn+32F/TLTi4cwhok8ZB+cWLY4HkSesM71g3MPv30T77hK2HPY7IbGgCpjK
iEwB6igozyZCbXlXXgASdDj1+VLksMdgC44Vhu8KwRnFIiAPXvbV3vEqac/fZIhd
lhIy1aBfrEYXHXtgRkfzSd/olShuglwvVcF46jcOd0hgTIJrGgEAByEcSvg4q8WP
KaKykI/JfmXf85tkt2kBQWKOVL9DF2LxHUEtzTGWt1Qn8pOQI65yhlkFq1IwAaQD
J17L7A/4BzgbZYSxJIoBCH+t2bvYjNaVMMCMMIiFaLye3+COAvcigzJD3mHggUUF
51GWhY1ezuEQdImcf3YBj4SPg4T4i1w0wD2nSsuz7Fy5tGAps9GLeW32dlSprAUB
8RPVi58G+vKWQVy1YU3XArsqwdM1uLabsFIoJh/UrG5RtCBndtERHC1Gf8xoJct3
RVIcm/IGVTxTilrOZ9Ps8p5DokSPGRxvLARGylaJ8vs50ujknYfyxxvlXfgfYCZD
euwKUE7KckesXPc7X6+yPkAUUZ2nfJF9yWX6+Fwpuw/cIzmTSzPdEIGW9CZO4pZe
dvHrq+es/fygwP5a83JDBlnPPsLfapEr0Uzg1kD4JzDWV/i5RKPp0RdSo9bhdKOb
0FcI5EJ2ReXxb4qSTTGi2JsC54ZILSmPoqMwc8EdWDIXd3/+1ZG2QtvY8D43Drwz
64a11s67zzw98JdtRvCX9D1j/mZ0kN1dZgbk7pfRN0hThb5Emj7O47fUl+pDZHYU
0qgDNvtV+sOclLIhhdHJ+F9SfRshD777E6MJziWbyz4WyG0y3Tqi0PcYy5vcRjFN
6GWP8uC3kOtvMAs1bfzqX++xA8xMajR8Xb/LRPXJG9RzaDzYpBhPHYomOU3QPNzj
ph8g3C7KwZX/HI6/91NpJntfORa0nNMJAmttHeU6srhU7+3qhhetpRMYbZRVQCch
h34aEpFAFjLxYD+NI/bt1VNicTrtssKQDe7UhBF1TVNlT4jGPpPB0qEfITLDUfFH
C118p3hTkkXAV5ZK0mDKuzLZvOGG3q+7m1IMHXvvu0A4qEh5lsMTgE96r5G8dep3
ONg6+xyOLZYZ6n/MB5+/+rMzTK8Ph3g7v39jf9c/kUPh6OyCJy/QZhuMuM52CeNz
EB86B0cRKBnsmaZVUwKB312xCC9PsuprPyOIVQk+S73+qBQno43K+5JoJ4UTJOIS
JspY5s5BxIETMRmgJVoj2RzF6hhIBPxn7c4ENVlRBd7nSVDURx1e2S0QM+GYfFe1
eabYLV1RPocVjFf8GhqWTskv7ibLq6mhbklDHnaQ9T0yg5P850nOq4SzQjFhW413
6Dpz5etIpTMOvytQZLzPFsYKlTEqVK2i3UCJX/KKp0xTHdW/+0qB+dINMWOlH4a6
vNnKwzzY8yvKQftAH1OZIKNshBCOU//KveCSW7odv4OXk0UI67Xv/5IqTFDONafh
9nVKWKSTC/t5JZ6O83s3rlN6fe5QXD0bpMpA5a6ILLlrlrMBQXq4VMn2t/1wKHdy
jazgkAfuXE6tISL+mVqe4Sa6xQYFzxc7ZTWa3IFpUiT41B59I/QeLWO2ETQ/S2j3
TXTGqnLscRx528UHOuMeUVLnZu3sk2Myq0HWU8a/yFPlgh5NVIfQ9xRHyZGufHP8
rxI8Ehe/2cE6IFxUt+giW984Avuivx8qpni9HLLZTtVeoI6A4VZoZEBONWWM1Grz
yUZ/ZGJDzf1oUDYjX0YeNFOJFlN6g7dkyx+9RNNNysbr8HkKFLaKuX2YmGD5SYUp
afxaySltvf98LOGnlZxrkZAL3/Hr2dNp6QwdAPZ3bFeXaoGQU2ihUVLHeGbxODHv
4Ym83xzV8sdkcQdnRriQlfAy7PSNoEEhsgqUSis93vl4E9vts8ZJNBITiomCfaiX
4lsqeea+81q7ndPxCJZbC+jcn/YQVuFZK7o3Uyh87WqGR1812j3wMxcc95XQtMFR
813h3gtmwepTWtV+2qHOG9EN/Hfz9zoCQ35ddhnNtlORWc9lEm7hW2+kKsHilXJK
1bbi3JBq3m9Eb1uhkt/GM9os43Y2Q3ew53tNH3M28kSIapzFf9huBHk8bcnwDFEC
3A+Zt/UR1Uz5ST3vOY/NOI0yB2MeDu3OIDJyuJcsE202XLmzLY5hC81XJku0Jid2
JgpbYMwWqsUGRxkuzyZPERX/5U42JHNtYh1Suc0AA9i0J1DA8DO0HUxPO/q6muYu
Eq66NA5AzW4gGhRebUxjogcN2/ytREkfaJqTv39Yoh/M9rkYu9pyy1p8DpSUBT6t
5GruckGu/okzHy7B4R7N8sBHC+/SmGkrUloRoSnK7Mr++NCOj2VHns8jum6Ke1wf
kFnbu4WmjJpBHrHFiC29qX6ULzcpFjmqprG2xSFwtWM63yw8TdZ8zNYw31e3DaLq
kY91Xm2HRDMCOMEsmGzDkjqwikjT6CKxedFmw61BVckgnwYIStDAl4xTfbJp8l7E
cyCquYUXHOhYDEywqHG2i7CfCKvxhOmoKFyzBnf0yiys+7PwoY3OwwMS9G2/ydLR
+9My+yTDVrX1KwwhxTmlih+7uKdCyPaMdCdshEdGwpkOP/e6C16ys/EXlemGSlyH
h8zG29Yu3+TzW6wJC+QH78WSMnm+Bx3vDE9dCxzFhykGF1u+tWwClJimRlx2W8rh
tP75fg4JfLwfOuQqlMcGt4u01jPgAYZZbMTVpzPLhWlozONlmWs0lykq3GUJjZyn
T2pEAiJtAUMQ7hZJs6bFPsX/s188tAbkEBTrIMS3vL9rNsgNsgbjCiyD5DNP+rsR
U19dsb79UD/hu1ndmzx23bblta7ZgGGFFpzGJfa6VQFoV89UBVcx7Yj7V2x6C/tY
rYQPzi/uyKVzJ0zp5GUKUtiR5CMZzBwddXkZ5SUFq26RfLkfKye15aH9htfrfWL6
o9QvOYXPWPitzDdA/4uifT22l15nrGeLayj9P8yiY+59FYz8aMJpjnZalRGvKbRz
hCnEfLaUt+bTEjrr7mIBgglBDv6YKnsTOCE9GQ1UyS9H5zvrrObxjAsRotn4WEcx
EPKRnINuKzSiCWmnZQNjIqZp/M1F/UeyCvGiBmgiEVC09ch0w+VYp16VXoiQFBOm
8JGS+wnFkL9BWciQeTg84m/c/wsgNLRyxi3fiTS8h5drVqE56899V05djhFsQFoi
DBKGVZEJMyI21Qr2smIr7bBaN2nm1Eve6UvWz38xz+7m7E3rMI5I04hAZQJcDUsK
zOBOJhSzZsk3e3/koL4SQq8ZQGpaEMU7vzLpjcUQuFSIEvyp/r6dXCku5ueDsTKN
cbQbai4wr0m7zhAvWalMk3HIXOlK+iXFLdRDxeM/N64dpAdQDvfsZKBUIsbs46Qq
z3hrRE7BsL7QCIUS0fZfGX5g/yL4oIltJKpheN1eBPSO8WXXM9MNPEWMQZ5oTzje
lFxOCyEGodmBzXijFpYeZSUwS4FPCGHg3qpv+OjK5cM1WO0IxZOK7FzIf0bKlDie
CJkchJlfuDUk++l1uivnJUaNCpwPcfl7CHZ9075lxJXRZKHWPsB89wwSo0MktBmZ
IZnAfhyH4y+6eAabfeVk9vUszmDbXBqISZWPRHS4RKkA9/OtQyfG6e4ARN89W/0h
m9q8WDTkPqbD5xIc9y7sD9s22KZ7D3BWBNa+3I4MH2Xx7gruXPlmnhQQl30IcYFr
0UivqUAYWkfPD4DizZtRy3Pzl3YY7eNSqcpnLuiW6VJOEEOEfFh3pbtgMFGd5lUu
fL9gxc6Q8Azu74iPc6uIO++Xp+KsTDqHatPwZn+yl5CJGXuRHtbMYCqb2jqiJRVV
LEM3EZg3NStlObQkgvPDYNbp2s402ccqamJK4vcNP2aGtLINMHE/pJOvLFRfqEX0
CWwYpembmgwNTyCzeP1gio/3wRkvXVssmLdP6VXTqY3dEJxtCUz7C5rNTBsjdkiV
/UBIpMBolw+5Y6dG/e9EDYYusPuqkVW/tzlrkafS12rdvuu67sOxkn/HJrDLueGd
454a1KKzhoyJbbwgqCJ276BIpgap8xBoAXRsu6+V2Somy5RTgz9l9EKNAg3xpyWc
ncwxQe36jSpf0lOkjBxS04ijtxlmlQYJrMLue/uAXKfv57k32luZ5GDM1i2b2m5y
gzPnUlfg6dXaVW12Sx1XZ8P4lUaOTDOTod8k2h6KHHWecl7ocUQMIZYcsEKyyCNZ
tmqSrzmeFO2xvrsCSDVRM537fjs8TLdukePQlCza1hz1ZE9bfYnOo+8OSeRUg//v
Ru4DdbRvZAHfO8yAUbEUeaXX61sceBMASlT8eL6DHOnkMZ6/1LzwHUqlkczkb6cT
auIoCx8VEpSLP3qZqXlTdQaaaSl6eaiwUtYpaT6uGQkm/9yZsIRqooi9sAfK+iUA
YPAY82oJod1Wg9G6f1nOv0ZNvjLn4znrIQrpSQYj4T1sRsINlADJk83I/ZBgs+eS
vt6Gz0RT44zADb1M9vDKm9GbYSUuiXaeg+5duLPA/O2tza8uEIA1czPtaRDCyFbV
Mw4pm21khzlthAXNukEMlAlXm83FrqtHNwp2TXlAV7qtBS91vrH+EoM1mm9NAUrD
tOPcpc7ovWGJfqdDqkLeE3vynuQafn6Y+uCJCMGL3h40X91KmQn6k45roYT8Yogi
JlIgWesuqCQZ2lfEFzeDPy8eM0DSerXWe8TO7yys8hk1POxg2VP07T6ZE9rgPTrl
q4v+SOH9HGjAAe/6UgXgy5B72UDKFQL8WQ6ZM+vm1hEhV1RcGTEmXoAwNFcsb+8B
r1Hjr1ikPj1tRzbMDxxWJ1VBn1ThPpScL0mVt1SZJBruq3KPyTuW+RUGN4LBDPHN
5RAzvCpKecUSOHKeo6L+EuTr0DAECzk235jqKylb0GgqVNCuH+fR58fqk06tDZXm
QrB9LrHKmiKLgcguxFgQ6SaGE5fNawVs7+Vu5SXWTV67ddT+bLbH3DT/5LqyHvrF
ui2T6xbYUs3mWUqbMjf+/t2wGymoyvw6SMxCt491lTHllk831qERNC+Fd5I3Q7MR
r9CdQmsoneQDryQ0P1oy6lN5t8ZVlpnyFgv5DP1s8yqHvHgr4PhZSiJjDEQ94N46
9U3aZfKMS3HVOFm0OcHw+11MJSnB1scgG90Ye6FkXAWQLB/h9oGlRK7AG93zqwjx
YeKe30QXY9AQzqW9lRrC/DGRGSDKXz6hAYSpPusAw9k2Mzyo3HIFRsn/k483RFzl
1h+/8wVwL+B4wTgZsqA5QZzoeTMKCPC1ScTzpazgQDtkpGbkuDs4j8qOJYZaoLCZ
Eu0iBDW0WThqTnkWhwvV4EpUNE6uViaZ1NXLAzFU4Bc4iRFKMpdDzwxxgcCn8EXI
kg1mm1iAy3QAGWh9jAoIX9YIneHykiQpPUbugdkoZEBGrql5CJ8lxWip6nkrxEV1
AqnaJQuhJgTgep4NVxKXcSh02sAEpZOuiyk04hBred1RzF3PuZ7aZc8T5HCGKVvw
UUVVaNjLNbFBis1V/QKjF3HmfYVjtFBw5/uQkveec4hv7Tuah3swY2TyTjL13EFo
EljqP6/oSTo0k2bCiS654iOUqqLTJnXkGHwQ5+FUkLNleGckBP77ZVdW6rj4cKIs
JxcQqaQF4c1SqEeAOd3Zurn/HsEwwrSvkgtyKSZS1n/VOXtc//df5/nZjC1fciml
U3ice8EJMD0nn+cZDhC9KHO+oAXQr4Pss0AJDklE6fzDLrQelkAFL/ymvspYPp+w
FB7Uza3AIRcwcOF7jgLYsqH/9IFCwiFHiqE6NOxnm9TsjCWSnBZHjCEVSxMZBVdU
Z4uQrbw6xmQczbeftRmV7pfRu8mq3uD/lRRpuR6CXF1OJvPF7jSOdGPmTspBgAvP
Hgdup2jIg5HRlNVDxakpHoJdo1svUgCaz0zuz+6oKPc/Yg8sCHBaDdARUCevOnEa
usZ05mtNb0QtgqJ3aWFjb8Cx7vDhzqwv+uhqAA9Sh3K0kUMWczwx7ky9eCMCwPGC
cCXQ/jq/GTtn32S8pna9nw74juURqtj21Yl/WKbiqlEYRRynoV0lML9Qe5IZT+xn
fr/a566W4JDp3guyFOZUpWdGIK+trzdol0RVN2ZtYEsngqhvugsmdpP+Hv4VWKLi
AMKcB85wsE3pQ92l9DEqTMhtoJE5MM2R7yua94gXY4XQowpAWZ+IgJNZyYC0zFTv
gyq4H9kcoo93B3IuoBEp8qZaRRAOv1P1pDYrcAx56vNpyjIydJToRpkSKXPIHnxj
P0ggWKfgc0LGDDqbU7l+iSc/fi0rseL3BXeLv6qve5hTyhGF6lbE7BMUZEdRSjcg
R8H5KHLxwkVcXWjwY3dcMxqeroa3vBlxDk7PUbHYzQsTXzIPWNC9unCY+/Frgv0u
pkR1lH6/0m2w4V52LNJZvT8FkZyU2xaAmqQh2Wy08b2+o34ZSN3ZeTUpGysZrj44
azaLqnEXnXyfRPg5PmbSmcaY1IgL0WQEPbRwJEM4jcjGAPkKlTDqUalcpejQ7n2e
Y7rc8QWo6fxu/cmpW2x5xTNiAEVWsZU0f8HZ2L6eFejhZ5KCmNPhZcO0GKqg/5Za
BUclE31bWTTQz9BAj8gxZsG/EnVH/te1M8DCA4pd9lZu92pqA/k5kTqdBdImUhtJ
aEwp5aEnQFC/SLEsxtN7YUO/IF6taUnVTPgoETFmOuCZi3T0fOFi/zXqcUDjqe/m
wBFVu7wTWmIcs9ziSOVzjUfIAcydfPbzbLuqHg0vwyrO0FNe4+hY8GgZiqMgg79c
EzjWac5mHeh15171A7Non7DdRTjHLvVrbR0jysMlvJ0lUf8RkQ7Nsk+SbyPqtToo
RRQVCv7xODnQblenx1mUMzvzaOah2RZ9NpDr2OftvDEDgwhq8ObkqCbkROscrf4A
W4LaO4Bs48ZwGQBUKfBK0G2k/JVCDfEXPcSTgYR9nUKduy400xYYOc2QD65GenwZ
yQqdv0dHWw9aETUltqlaLmhs+ei/9vZmaciizfUIiOQ6yRzprmWjI3XxH7ziNQOp
DVMLRm6D2E4zQU5Iwl+n7+tIabPzu3rl0KKR1wP1VFPm3C0J5Dn+mc+2RrPmidUe
+E4BrTIAZZeFAToVUeQzG/Mm/dgQPZ6Iy47jYZXBykZqgnx9TrlaGksAPr3W1HWP
T5eouFzbSmxYZlvUQY7Qessdj+ZqdRyAo/CXl9KmBCO8R5aExR1cfWBC5Q69ZePi
3XJduu7QdxX/W7xL9veX0umPvBiBMYy6VwzqD8RJgaskHQZeUCVYp4WXxcM3BTgR
BF9NOGLuWHgOYUor4nTJx/8uKVnZRW4MRXTCje6lO1N313LY1ppdcSBP/5T8dc3k
hbUXIA2qD91MywxhNNtxuhiy/5oBZvtoc4FYxt5FK0F9TTMmK6xo2ajqGMvSW1JJ
8iCuErqiICGsTZTKvvQ53DUV3q39Zz5Ghbl0R+BU3ReaCJzJsIq3+FLGbYMASR9f
aRmuU2xAnNAcBBId9paK1kw0P+MfJfs8o/A6WO9D3JXnAcd9PB3TNp6GsjJdSZsF
2/RLnhCipGUO9iCf/QbBYkSBeLT/7fQL/zTwSITFOHM3ok8Ka/jocKynX3z6D7i9
m+a80Cs1g+cbsOEc6nnme8oPHlIYZD6zBahMkgQ127TAnrEFpjia/xr6IBb2/zqy
dxXWqsyQy1bXdM2Y2CI0cYuExZAHNkd93+J+WGDnR/Gr2CHdzN2aogIn4rSnupaY
2QRu6Vl7CK1SUtfYFVj/2NMBIQEaIeU4sKIBNOEqRs+Ps8cFy4n2RuublYaPSWmU
iZ6hu15bDV9Rbt40jJUgKUNkPgHf/1E/5DWW6L2WVoGyGFwdBx3IgtBdGofAOu+Q
YRXv1cOe9Bt1ZFScBgeko8j/TcZ4xoP69+lUeyFAk+V3BSY7ROiFB2wAzr8+86ws
N+dSElzGegcSnXdcss+h/df6vB/duAbWvgUcO4jsuDLLvpQQWMpDRT85Ehq8BiiH
Gw3+fJOdXSHgGlqVhitQZBkfA4lCmZo/poyiWuLxz8hq5kNYES8Uo5VMMLSVhbGw
3IUxHXfjfRxxRgZc5iemC3eQlEVL5zvIdLnIRk4picIBVuDavZ+I9ZTyjQeGEb6t
wZJAheXMcKqT+P5Skc1mdeHAycSqpKXREKAipNiRAtzuamrbmfkJ54l4BZjD1hYB
1o+HPkM8MF1RyGtp+GBxU+2jHaQm8cn+86lQt3ORYHXSgp9MBOhys49eNFQZOBY/
2XcZB2P8i6b2+gQVdadE+x3eCm/6G3GB8qGM/1xgQF25hBnHGjvsA6rkPp0O1ldV
KrNFN+ydhf8QK9tn1QMiDi1oa0dN2hZjvDEnzi4/8cKYWOCM9NbQW1JGWmbj6faz
ZaWCJNj9w/qBlzgr0YE5VL29DrITDri9WovPpdQUWCjnicuzx2OBs/p1oBJ3WfHP
Yrb9MQRVrMd+HLGsy9EcPsI6KwxAkI6onBRrJfKzk6iaEAFKpHTBqO4E6bKIiE1m
RKU5vZGXSjs4ZnfLAwueleI9tzCVhCBVul//tZj2BG91IsoXSeAhDTyjak8SpspH
97B5w5FZbbTz8QcqLT4OlBEQOEX6GafQtHnm6aOBcMTM12i1jfwtJpzwrgcStE7R
D+mB7Ym6Hs3Dp3Upwiovme78s7/UkNZeqZmczpAzFU1iiWPFMZGzpaDbwEOXLiYS
IZ13O1CAbIEKPrIAEqgULX8b+wzp49j/Seg6IGl0cAxn2lFxOZWwbjuqLsjTjcii
cdLWdEQCTiUe06JmzyzXn4uNThFwsuKnKaa4t9wZK9OxcxN1jBpgE9IuDkbzJ0n2
geEVvGFka1hNtq7K/1ohwoTRZP2BLP4yuREfvy3MN3DmSw6z9+KQctJusE9AaxqM
M9ErjqKBDhUFiF9+VfLY8SX4KejQ93DQn+N25VvbNc9op2kTLoRtHiK7BmF0lVLQ
Rib76fVuJ9vMjnFGuJiyt37Xmmzp6KcdheJgQTZOiFMpqa2fCzNpmNx2JrQz+32P
uY24jxZ4KY+SYvNsw0EpFYlFlGZ/wgYEd0IC+knZeNPkkFrnH6V5tXdk5Dk7ns44
jdR7ZfyT06Piq8mvHjV9x6/s3GxEU6D0+P7AG9WoMTjHzvlRQb8eMoAAW101Yoom
VaTd2RPXnGQsTh/jxqzJqURlVN2ZdCFz+ecOWTWobr8pySCLSmI0e1x1cXNZdS2m
2DGpi9opbTfVpZ2ByoLf/tUdkmRp2zts6CWICX/bJ/tOir8B9b7fhVltXFnazJ+l
mg7WPV28pqgYs5WviyCFGphxJJ5c8ZPLzsFd9ltsXWBcFKIIPJtPP4wn6IaAC8yc
RM0zMnZ5w9bgC05pJj25JK8W3cnbthoL+gRZzCpvnIuKbtD+leWhBBY6Nd2HZFfw
YnLCQfZ1fWc+f5WtFQUMLwJbGcBm2RuL0wTgDVhp3PCUUYSEd6OEwSaK8Mx1OpgW
oiuZxOFZ7QK4UFsLQru7DVWpPGXP5xamLLxfRSiNMXeP4eXVJZGUnp0sr4rhj2hi
KBB9K2ZGYAslQ1L0jjW+ymbB4KM4WiVX6jutNPyq2msd/SBtqELGJ1ErEwsF31fW
6aR0VLePpH1vc/qn39l5YDdyZVojK0KrQ9MGMw244jyTQyk2AhaVLGPO0GIJtxFE
V8vQH1qkeVJwLkFqu8OtqkUXo5Fb3f45kixKXebLRjrNrVlLKETfkHYB19REEWcQ
XIo3QWQHZsrisRpZcyW+LiUqx4D9oreZfsW78rprnrmj2fSsAHxpMqvbwTnGl1pB
70IPlQLKLO0zvAO4iwNKqu6z3JlwinPA+9DqMg0m/ZrNqf4kVqUEI6vbxeCuMQzB
sCrxb2Wfgv/saggNkNOQQSlpZRq3vp7ozEhqLbW6IEmt7AWCmkPu7TjDmH/FsOGK
XApCA3iiEOR3sWFqrEkfOJ7VtChwaasvrZKlN9C0EmvMJfR9biX63wcXPO7PnouR
cSHmuCaX5i7LJIdmOSs6ZsBZx5PoX0GZuri3GjOfFPi//FkvIvrqThNkGPnYMwxo
YMAxtxWBF2ywBfLQnL4UnF0tWi5Hw5k/iki0Q4HhnOA05M1edXdhxpEb3CI60u4p
uo497H7GadZM7FpgsK4CXGdMBHyITcIzQoJZJICKhfLW4soJAeAK3cu+mZgTwwIt
wVc0WI8BWB8Kvr1TurANy5ipOABdEaDEZBOP2X8dqpeniCnUFLil/CffAmlMCdXT
S7Zx8O9l0P+f8e0DQgpHVtOpeY52TA8oTKeyT+XPyh9cN4xBwUifU0wo6BTnmzwx
v404/gsPoKWFAAVUoBE053gSit9EQyzG4NSkRWIfVdBTHvamVykkBJMZrzT6gc0B
xIeTjL8XsZ2SjVIlmfWjUZs8yLVIkxTXRLmI/inv2qxRNWjO3fHiyDJ7kdNrFmL+
UAjDidmVASw3lCMP1xrEq0/BDbHwWNSHwbzqvkTgQtKA6BYFmqaRi9t7BZf1sTxq
mEQVaJaFYWKpJNew+IY0xwCUPziJ2m7QQ7ravDNOUqnXWLU3MmlTzbgUlY5VvXgn
/d6IcBuxAR2oTwz0JZwxL9MpqfjhnBgSOO+KOuht/VnuSWbcKy8JN5DT26Nmxbw9
KaJVnHDKA229M1/HZlV5gxL6KgEz56h1vxYm+Hn+ZSxBuRjCT4XoJQAO/k8Y60ew
rkSEmjOioO2ySo2pk/hccvN2Fs9brCkCWUY4XQrhAlqFogFa46wjuDBuYTRPcFfz
ZjHm0pu8yijUXHhAfXssBN2uMz0yW4OveCJ7spmjoZKFOb/+CLVSKl0RkhbXMB7Y
aG0Iyy/hDJeHZrUA1RyBvkEx7UDEm0wkZU1t15yE9ts+Y8JxoTApOTy/AUvyCOfg
eA0sHtoPrKx4chKqmmAyBkKkGaEDiuQjr8A7+aQGTanwKd4gcSQ6CEUR70eLG09L
MEtoA+fx4dIlZFiWXGH/uDIr9PFQTj/sBi7/z6hHq9Oie+Uyld9g88M2MKLWFbWV
fdPi5GejxfGrAGdV673nS2Ap4j16REsn8Szh/ncLUgQUOypbZXZVRMXrdHpTWEAS
xDn5Amm3A46Ui8P1nT3pYinOLW+DWClciD9cSba8uNsosUWhDvt5GTdHF3niYH6h
G3v1lFY1NGVz8ncxeVBrYyQKPR7visB5GHJJrXxDE3HQuhIrwyCejij0Qe+p5Dhi
oy9fLT0n/j306RneEm+7t+e+3SNCrIO+5gJUSzp2XspKIKTVj89hIfbg5jdRi26v
uPzU2FAHfp/6HsgAz5ZdEhhgR/cgA8Q29TcRJYm/F1tUphnia8r7WC97hTJlk5Ew
IBSKYk0TsKmDq5VZJz1HFoMwZ+Tblgk865dIYpXrpgnfv0VdbSlWZIUUTH2bZdIC
4zirNP+XSCkJUUpqV/odT0c7pkoEUs+UtcqvCHvIB6jKbB4vXGGOS9RZIj75ZrN0
HS4x+sR9AGjsqeAfaqEbVSq1f6a8OCK74gqfnoXMiRrKLmnCck5xbbUbOu/uI3kQ
odgXzkxTQLbHNf8/7rvrlD+KWEO2rgfrRmauNPUpfN4ZiNAL/zHGHnFvKHoJLPSo
Rv5dS9/FfTIuSteGKSZH+zmaxJhLTE/FTPQfjn9+73qCOnnUJz7Lc0MCpwWoCEVR
4eBMNfr8eNBB68DIKa2f6PDJuaNBLp/vEqEJ7/PEUmtVLGJfqw0tyeXKDKhR4XYH
SCettHTIbUjs9ExK7vTKoB2kPKbpcz+asAq5eSYGozkJB8ISVRd0PsUWsjp7yDI4
qAAsFA29ZPDbpzn7ZM8/jEMTBtall8ULC2ERv+zyBYJUBr2zXGFpNN7v3lZBxOD/
NvB6PKgee7H0jouKb4w1ylSJAxaS7UBxK2fpMOaLgbcjE8F4szdamiVlURx39uqa
UxSPxDAIbFXBa+fuViZuo5/JlKdLrc1bWtPmt1khbksES6lZIGSoqE6g3MWQFt+G
j6tJPjnb5aJqVT6+4ZzgomfZ5OzgV0Pv7lhxsRkC+pLRiT506STWy2yn1AAY6lC0
63p94OqdRinvI/QxBGcDot7IABwPx1csVy+n95NjNBEA8NN5B9dmbqGp1W1yf5S/
lAgbpQAHIpkK6E+mds9izGz1c62rn8TGw1XM7yNdzJKGHPAlcxBQ/kyooBhV69X7
Qk8gC6gCScpfUdbmd/68egh78lRJVsF0hh6TuSB+6V5kusuhdyKPn5RiWe9p4FDl
ZJuspU/DhQmcIvE+kGcAwXiDOXvttOETdQoVQmB4T7oBGHq4Bw3xIU4hPutYOcsW
1y596xH3LtISrmh50H06xTt0y4148SrOOF/ssHYiUd2noBuglNo4BglJMAlTCbHu
FtvONvBKvT77iBORx7NJHq9AJGqUP9VyvKbEc627kdZ7xDU9tcsPB+m3VQkcEtWG
O9gvbdgto89gLQGWOMHNyGsHzlW9FmCuXtZKfSVlq3NzdGazCylGf4OFgfzqfcbo
+b2sP8rc3gNv9zb/fI1CNYsGSPZJz6wyEygY2fXK4j0M6XLUvo6hTduSAMH32/X5
eXfQlLb/gfXj79jAQaUkEbF9Ck7QtJUHyNXRxlmLx5r5q7EtC2mv0FGfyRaBX8VW
inPhZxfylzN/x8PXnDeVzxF0SqZqj/5O5KBbhRV7V5emHDQWa20/ki5aQlWERwKO
B7l4eBv3M+115yO1h8COTUKMBNNgZh+n66bMU/NuVRgeuppJoMhh5eeHykIMvIs1
Bf6/dpZzoTtGSI0iSFP5eHdqJOUxJKmXG23E3uF6OhJi8jWDaxZxhggjjfnEd7XM
OEAkLljO+xrKLz/7279JhNVCxFiOWFlSOIAHYx+KzkIu4Hflx1m84NSAbQ+rZk20
UkGDlM9uTzTLlcfCtVypSwmio1Mim//jY43zUIFsgEcaW2N+H/VQVg9PJD0H+eLP
nI06iLS7Ocdmyl+B2gwJAYDQ+0CKhJFtLw52jC5X3Eiv0+rrWh7pQ+I1jWj0SnWz
S12jRnrWCHIovVO9l8S120gNtU3mn9OBCS+683mOFLP0JggCfqCBPt5PPC6MRyYJ
RtLDx+okfkkqW4MCGaHRniwpbcKqUhQtXRZmAo/b/SEHSKFIF2MtAPUiqwef586Q
9HgVn7YHsY381dm0+q5LDsc6FmFBDS6M8v0WqWqR4gOrByU7Zm/IRRpVM8DZZ+RO
JkKUMsXc9tI/KItLwsumtBN671ff1zy9KEsL6N8t4xh/swlluhZiI1q4+ksXzd0Q
6yJoWu4SGdaqkQI6K1SeIm4P+lwd3TfhjZNqGEK1APpA/gk48M4AXLd8G6+8DZrd
hjmM9XuQmNLFUgKQYzU4S/GKOSplNJSeYcotKrWZUlV6OFh27jq3pppK4ECRf4Na
8WIlV9JHAv9z6VAr0nsreWqDKoZw1gTUtSNIfjivctW98FmHDwpsC32fx2ELP+PA
ydIp1kknz2iRRlBwEux+VP2LhImMjOa6beC77fHUCNVVaf71E6+BfSJ3ruoWIU8x
DOwizhR4UY9s/bkzxYqQM7UJJFPfsTBdpDdgX+2EsHbCmT/LYIpuzsvRX9o7yGpu
v2aLX5rV+ddyjedrO97RDtbFbgLMsw084O1WPqWkzebKQ3WSUjrh0f0KsJ5lejU1
DN/St8qZUULHQY77z4odm9UQi1GbJhqt5y3EvqiQdBbqiMJ8mFQglhiqK42KjfU3
WpiQq1LOFqEIMNrAA7jDreXRS/nNSMUTm/EWSf7CXq7o12MYPXe8uzpOlHkckLd0
FsuF/QRycnV5DLOFOTg6a7k2FwIOuw2CAwd8p9jSfx2dRKDFuaERKCanJlYEzuU1
2y5ZBXSqjNJorgfboj8mDx8WDp9hKvg2WReWoUJDkWzlrWe+ZKN9lw4IO72D6LcI
kjl59iDTIXWJhZIGGDOMS/wVaNRZzRT4Q4KLatLGveZuuSq/xxD7A0al8AYwOypT
IfZYnegjadPm5w5qbPCZNwk5wQ8xnuuCXtmJSEs55NvQzFT+z+0jg0QRE7IeY9U/
Hj5EM/vIzsD4P83ZyKlBBCIuhmf4VXBX9h7l6RuSnnmZpwrUvnpjY9x5FVEa2S3x
tPwgnqN2crv3c1UJWMgUjX4gTsXvW/NJKOmVaQOUI6CwMgRCnu2aWnd4Izxlwqfb
Htfc30nURi+yWk9el+QF9GlO1l89CVl0BmzMJ5CfB8qWJeJOBx0nW0iGB3/oWomP
rsVreP4Uq1Z4UCDexYnOzhtIt7gMeelsdDBcjitoeRuRV/uGTg8McYtQDzhxpsSh
VBhmWWtzYBQyVLcF1NiswbjkivSHe4K01PFwPg+FwaCNYmYhc3tM4T/H8QIxIMiu
6mZrvOAXvjnmgi20P6Ffl0hIFn1X/l1GTFDXZA5hdEulqASGdYbJuV+k5U2MHHGY
DILRfHMfp9hBplXiL8Rt2l5Lh37yHZId3iGMpuqldTO8QaNKtFEL8WvCr9exRgo/
ntfThc2Cceh2jMvqIZjk7WZBfxLTO51o/ogMQmHLJfAjUglCYMFTc0RzstWfCx10
B9y/c4U/2gV4B4PMUvkhs5nkWBwYY/6LV2yRSb0/H9ZgiipZptWo3yLXXwgD8AM3
Onocwh60TCkMeiBJrcHtfoQqgZkDpu/AErs04BwllAxSzG/6bEH/NVtsPcYmswpE
pxUKgoBL41+ae97jKqI5p79o3Su2pNPrqwKemJdDV+9EOPYMb/Whs+ZH9CkTh1v2
1FCmfVe/LSIyxewEzPi0UjITEJfG7q9FNHzPRJuRT++c/vWByXwOqv2UYR7Ckrcm
MPVaWTWn7fG5sPYYPtL9RUpOLCBPYFEuZ5BKGGjzOd3FY755U3AoZdvITzbIEVfm
CZG35ujjHN7Sw8JSnflGLqW21Osh39Z7MtmUclHvXKgeJdxbsB+Xz4VjVjEfNYvL
jLrgdtvD1N9uHUrruJ3J646N439mB4oaniAnLooRu80Gmzf3j3K+2ueuY0NoIZjX
byKKAsNqddzCNMzd/1JPXU0k7tNZfsgo9S9+cyeDv+A329TmL4pi1PJHfwPKdF43
BTLtGRWs5cMJMd1a/QagRq/ZAvPlfO/LSH7Npi7YrT2Adq7MTzkYc4UqBaHrzYTz
psCqy/QUyrQRhIKMuREGHLVFzzqTIbKsycuMogmhsEZT68A1DeUQ51Ix28l1iGAn
R9SXcq7gttEgEulWktbDLRF3dNNhlU95taeVS8poRLhojyT3qU4MThUGj6BcDwX9
lQJlO54TO0l7E9bEnERWi/GQro9SCXuhnqnwbeUil2GfbnqlBsIj0YNzdZdUI+eQ
VnXvZkoVYTpS6yXaI+zhiFXwyGly3L8kRv9lJu63dTccH+L17IC7tuwuRSz9d0eb
5627uMXereZyLvXAS6l4ilhG8a8Q6v4/33tvtWbpmuxb/d+256VZ4RG446g2Grt6
EkOTZXtbrRcZygQwbw+n5wsJ1y9mqsdpXcKefy/h9RarEi6bjuzzQt3i0I/jkDNJ
/6n6QzTZxOMoI6MidALPVNtrjuSzv73EkUc+GlvNzf/RokU9chzj0O6a/AvkMX+V
uD4yhevxBjxp1u8czGDLDV3v2b2hs4fIap0rE+H20/P2nxsLHX6QqCbWYNzxmPQr
jwZBdqeezQ+pdDLMJ0PeQtST9+ja2FNIS8vdA3GGStmPu0z+NV4JMg6LKoksTyGy
Jsu1zkCP3FnzmX0q5pbzbeDRmZmm1+ufp/HeGT3YvyMftSz7hUbUVmNcGm4POiTe
wIeMdHcbzfyyQiKRq/5K4WgaLrAzXDZNz4iBB33V/44k0F2JD7Bw3cV+gtkttMdv
8JJLN2oZkI/MkZoWaaxiKtHXJCtOTSj7C3ganCBloR50FuFD5jynRLuX2xMK86KN
jMVH5xgEGlobfCygjHpzXm1RyhNwdwKIK4bJDLYr6ZD0GeTmi9kLHDFZoH+mx8Jj
CN6qB/uwpc6PefvnAKMis9yFN/I9vN7cC2H1zvlpgKepzunS+tq9WLVrOzLIKWSa
vyLSAXegBPERicFS+LncMfDC2qDlcP3oqa++EyMdvUGnfHZWei/B39Ts/cxjg22H
5xYf2VK1hB5F5Z9kqCIhCPcb/PNN25U5rugM1KlSUUMQ7TKqdAeeGQVeDpsKHIf0
0WYQOyE4z+oPkSDdm8jTfT9GaKN6ueJp/p/bdjeJBW9i1b+VAyNx+waq28Urx6rw
RYQc5xr8AMsd0idChK214kixDEkAfwWnEAQSuPOZ+3RgQSi514EmQ4ZECTxgF1YI
0T3ylfM4BthCfmJkzAQtrjF6PwPJy30l9s6eMrFPOvnIfraxSnk9M1nysWehUrES
TqYObMOMc10Jp3qlNVw+xpxHy6oAQhXhWwVMBpBCykJ8Qf37a3tMrKaxl1qzq/I5
d9/Bmoib9y6T6R3tqvfzshOMHi2kE92iqXYM+MfOa00sk7/IyyUZq7oh2ADw/1V/
lfiKz5xSlySLGqb64XDnqA/aqyhmv4lkCIfgOE3xa7+2PfFOlh/LPai2BeRsP+hE
DNluuKdimJ2lVxotOcbFNsDVGDkeHp95ex41LwOEliGe18KQI1TzgKjntHwGmrtc
pc0jPkWDw4SOQjDJC95239+7Mzkr15NZV0mcukoAtQRwYkY267vWoiXy3cnJI/g1
ffT5eOX+MoslCnpxWAisyh0DFVJqO5Y8TIJVhBeyYYyyG4dMGZyPZwJ3GmphgpBu
qSQrgbv2WRDrJultZgEKqsU/pfT8TrvHxuXFWMkrmfwqDT8zxQjDBVtTsj3DOxGv
RMerO0wYzNQbpgJueqgcLBLJdau7FcnmoUaKbw92xkV6777wUWXQxMJkWwYR0c2e
YzMl6GnKemym/xMYglvc9PdCUwMS5uFOlwtwhJ+Tbwx0dZ3Y+sDkfnNT4aTjHbDr
xhxOHeACJaFSjPROFtLpcxOvv4tKpT/fCpUQCB8VuPKWA0ij61r3/qelFxhSku2N
e25p58mEo7FWzYl2ukh3pHgvWhuVJiEkdXZaX2OyGFH8Ij+TbhhFHX44KfotJF48
c11q4wsxZZtMtLtkIL3iXKMtnkRXHWYXHScX7koAF0PzRcfjNrhq1vVHFhy0CJeb
AqKiemL5WRsB2rXImKifdlpGZdOU9AyefVbgxjv1v2gd8Ifej1g3vf9l4SUix3ZX
aaP7EIVFMopDFm+k5h3f6217zS6WIZkteoSUPIt0PIP0wc9/AkCiivAIYvd/rZe0
Mx1g83KOp73LNW2hz58Y+TiDoZpgnCuD4aRn80Uzcu4qCyq4HHEKQQfEDcJ5EwCw
lPgRkAKIkFfd4oOQtv3SNiqWrXkzdQVfggOqqd4N3/QiuPTxEWIIv7Hd1pcuyNXt
Xoi7oVswQa6mME9S3s1B2s1itXXi33jra47QZ5NNTWMQT9sMXkp5Qa8rOfxIw6L3
IWx8W3bcBvLy3YR93EosHPEYZXl006oK/91UWYsu2llbKkgzUuQm4HUEx9BfPPKz
yjxiRE8TMDPYKqD8gwPjt96fnk7hYsjv6HFf4scCOkOOKCy6iojpUJEEUzF8t7oH
nBDboa6U7GBGMi54sIzDC2EUu2tWybqXs9b8zkb7LVtKfja2INzckAwog3LtrNYy
xgzxtj2zDV71EmVh3XT/G0f8ssOH7QtPvMHnC1cc6QtQTmkvHqwAROTDK9Z3ehOB
e+BIro6+C9uXsN73w6ES7dXcazKEW03xxWIWs6L6xs1itnA1wS/xcbN/x9MgLYeb
ODyss93jQEGMEPnxZXexCp34fx/HufFdeLBQ9w6a/4eruAjB9eGVEwxBDTyeP80N
qpEfd5FN3KGF9DQHBwAaEfFWhUxCdRCM4gyNlb5/8mjZBXRlgWqbx9Zrc6UDJo2+
RaFWb5aZv9/egZVtUYxFU01CaI4FluY0BlhxDab4RFhh1JtedYX+ZukqZsLfDrwj
XdNVb0lss7w7BD9+uBVjGd6CA8/3ybGdQ+a9z3TVh909B/R8vfuRWWTCjAbG8akV
1uSDsIf/pMhjHaBWbvUUjuhmfmLo5C8fPhNv9ZRh757O69Rhm7Esrvl2BEkOOple
xXK9XuQ9BhrYnWGd+8AZIelGW+rwvROEtMsgJ4WI8OnlXiunGxaGvkmlQUTLxJFF
eVQEZxmYvoqyJfzBSaQ2nt/vy6nxm0P/BJGKAZVnr3uRQ++Gn58YnynDZDViDxtj
GX3D4u2TRi4K2JDmuwIHPDPz9+m++SSdEzpJs36XOnCuiwNxSZYMwiJEl+RDfzmY
3xfidTYCR21oa7fA/Rv3Jb5kZxFotRksHPdiLoNCCpxNvccn+k9hPS13TQ8hPi3U
SCuF7a9oi2TH2XyNz1pGFZ9B2QJ50f+fD7KMzS3/XHRPMQ2VLGxcLw5NvnofNHJ0
vSpYi+MIUyRVSsI9M3M6rMtmma5unuos0HKuqX4AY9Rv8MCIaPmsNDlzimoJMk0r
0/ZaNTf5uVevCfF+8+imfUArKAZ8xqt0xOtHqLwFLSwurWMlX6O2pLsxe0PFUX6I
/3ZGsEKXRulLlzKilcnNf6ShnywO+OZPPOI0PZp96TVJ4EPZZcIFVqBOFNe0uuBs
LZakd8RMsrO/1dqgVdJ0oncXsYY5CEK9067uzYbSPXFjS1TPB8Q97CUVcML7QwII
IKzj4zZixW1CVEPldiTvk76k/5OtCebzq/wItRpBVU94+nGTr1LHClxxmP4VFatT
2UFQlNxTzr8joxj40OoEfZ9M774YUp03IWPwp75Lw1E3iDLQPgLZKpTPzQUwrWS0
jHPlPtwwkASZZYT5adq+iDukbdzzrkUmpYH1ttKt8QDabAyho++kCpl1uEizwjZf
kepEGuaOZX61ibmranbiSOcHWNO3lxnybI9AEvB7HBw2TmED5vbtoEmEXKcxuvyr
5z3PElSg2YCpDIaYiUHb4aTHgsIanBuAJ9r0uF5tM4uxe6NoP17zkMBX8mLR24m6
cXR4puHGBhca8Q0+tTT7EuA9o1tm3diDTzndSDpJ/82RWHRUPHhTrPnpqldchxwV
Vfd1qWQ7cygqAXRQGdzoDHD6pLthRpNSwlnnTpXEwB1T/yZynOzCx9Gumls6sAYD
9x8V22rT3vtBZhlZQ6NGO+/elsDR5G5Hzd7qXas2E3hWVKGjJMXzrEKaN+LqbpGE
hvJzE418l0SPWdWg/h3XhNpfWSs8H72VjiZ1PDIYref946bFL+SgDchCC7rV7VBI
MdQFdC4/zNKNvNSfnbK12qlBo/nI9XsYKT29liu4ArtqTbBJnWSaNjKa5LIFNcMb
i977t3lNYfiosE+qFeGIShFJ8lmixUo8KJ+6bS/FOI7nt4a+2kgnB8TNyw2OiuiO
QeGeM5SB9wE0/I2IAYmYLMJjDu287NddgXpvv7opHDph0ja6hEufST1U3cJ6XY0O
0oMln8MtzSWJg48dxNItF23eJXugbfx09U83Zp4FKIqveY+OcDThMrm97XFVwZXh
CtdMOCg8ZD8VwT1O26o2XXmlLU+IKZ0OiiIINsosPigAFPHDQn4ZQ98NmWkth92j
E33Qecn+rI8vGtjk9EJpqg4Vvmu5OQfH5jH7lj4HgIAIJd+/5uyVnLu/6FV3gB7/
cbfxwDBry1rcb+w0qx1AU6drQGXhwzY992qT9t5S9UyO+5q13Wa4um8pk0NOsdWB
UGUaSpCeOQo3kmcAHy0YaZTzgp5BMHFYB/Da9lOlqXKJ6F9YW5jjX1nAYx3zPJE9
lY7ElvnjnG3Nj0O96lK5ubOssSX9B69JD5I5Hl9dXkfMIKZwkVXhWmmBFIvANOMT
y8NcfGuujGPYj0q8Yqnps1P/jTpc9aSClfm4iTykggcCU26KI5V/Z3vPLKKVNCrC
j0G4+v4ZYTIS5xfW0zywjxRuz4BCsHSPPMR550u3LTTEm+BhFfTqlrGWsFJ1Oo8p
nVnhodDHLT5LvpJBloR6hvBK1UqwNvDT9hyMnadSX9d6IroODaqjDRZQfqYPiGUn
7glVC+GfeZjNdl3CtRXirDsrk/lGawgwOVqx2BZCer9Kcgs7mF2XIw7ZPNY6rcp4
HvITdnnjmFZ50eH0IMozn20gv7mDeqldqfMyTsY+27fqZC/rLdkD72BBI5rTUKNA
V1Ase83VhiZ6YJyRUZwa/+Tp2ytRPRjxMogjs5oAJU0Pwmz/00aE9EzxF2SZDM0Q
9gfeiCIAHJ/IkeKXDO0an13tPxPb9mcfTEOeRyd7y3jL97iOxKPLfWPMMIgZRuWk
oX27hoaijGhCgZZmT+OV2/UpV1ORgL1BYswON9FW3V/gi/Rv4R52Q5VaP3fsS0yN
YcDf9IPmZAHiYQincquGFBAQEh4EPMVqqXMuHHJgiNtkmjc78PtgqAsZVwrGwRTJ
epklQnTBmwun0zMqS89coC4X2wWdYcwmujfIh22/+sg6KcBoDbwN/6hI5fcrieNo
V2cqjraFhsUzNX+TG4P2OOVj665ihNQAB6yO+bOXBvrbtZD2A5Hs3yLZLV3St+EV
UwPXlFnUHJ5HK5qz+MfVBc3AAYnQJYBzS/6RrqjdS1aAl2PMRER1YLSMXRDU6ydo
PazDR9IT3FUDYdHtZYFh65PCFUG5csvDR2MuWtJCkrwrcBkLmcBbc2ydy566xT7Q
r1XZ2FRn/0Z/8U77rDCj89OQlUg2RCdPwpG77E6WjJ6aRRWTKu3O0QedD7cgGu8Z
zejcP8SGPCexUQaN9Ppcbe8/3iGE9Y2IyYfpkTD4X5k8rLu050fWB3d5ts7cyXdl
wFQun+0qhKzb3N3FTJPvMM9O0OUs7IHtmuFNg8PhWQGwEoCVRXX4/ARnCUhjEvbM
IdCoY9MkHmetMzY0UJ+nNWzdUXcupAGSIzOM1CmtVGx3ljfJqBDCKg0s2nJvQkz6
l11C941kC+n+rNoCJD9wGonl09s/myoM/GV85q8A7TmGx8EtmR3O517guoCubuaf
B5ahOdrlT8WoTrN9seD+ZKyw8g5Jn64eMxa9L3hxkBvyzlQDgseUKB6CPqj5QNYY
QOfhilrye4uQ3+ecWyZHAp28l7vXnuyvXRH22gHO3fajKpYYgg4MZDV6Z/JGDZYI
Ej2M1oktB1VZ2pq8vg5KC68AETvCUwtqD+/nbXwaIsWDlHJEnRdi8k+qJw2HCYxB
FuW+4Zesos19fjhb2BUu5bPq8gavW5hPu+oJui3gIbeqqxDLcvC6RsGp9M+mAF7f
qYCUrpLvhC0gxgH3Nd3XrdiQdXovPpd9g/V6M7pGhyWeDmlhXoljA3Ea9QZUE7MW
6+ZiRbDgmxLN4AY/37vozLB4EejSwWxsCfbQHW3s06c34J6VSShlg7uF+JuqGt4s
DMLSJRi1qDfNI5gVfQrPbmihdhFsCFaUBCkn0d7YVaqWZJ81mh9TCViUxCA3QEf1
wdOTWrgoZYMRAr5VFoR+rkrrWiI3XkI3Ns6o5HiUsdaw22YLCBzJVdY7x5/VXnZj
q5E9Die8rt0fAeLBjzTm7vgI7o7wlExT6fidMRtRaujQhKntpo8kDgBlrahhojRT
N7hsMIU6oCybpdkcRDT7gZ3g7wpBqGU1JLzUtn3K67ReLBQORN4N7/CZorsV1DS7
P2CSFTMpQb9snVonUAAHXBtEwOxlQBjGRMGRv1zBwk+2OVRGJZa49MjX2gnNWUKG
bQLAfA5KUv98/rxVPjlWSihl7eGQwovIWXKyH5cnd8FzuPt/3VGeKGBjNKsZ7isw
Ke7n/xtB3rr7tgNHV0CoW+v9eD16NZty15oiDX30k17qxj1edX1OHmnYYWibtIqk
HH/mAqP4BcDbgLICibR3OHXzMqBLAICVBhXuzLkXGOS5fHpS7rkYx19E2m/pJ77y
VdTq4bP6t3C42XhJRhsoF25C8n8FpX86uKjsadEw7MyA8lfUVoLu736EggbzKzGD
M/KVkJgoPqhv0jS1TePsDwXs2cXw2kEE7/OLEtsNiRITaFror2x2AJdnsSbjjXRo
BuH///LojTDShLia60rCoXLpfi3xARDp0HuXaKiFe5WSqFtYvdpCqXAP9GS7r9wy
E6RWzGcUGmiV9X9Exmx1NRRwHW4nEo0+DKFkbPrf3gB3j/T0OEyHhy0jNhSXB4lw
Met1FlrVTucfjy+CqcmMjb49iTt9XVQ/SCxCrdb4JPMqjNEtJRR0n3INXIrhGTpk
hv6po6oE6vL9AfIetgqd6wpnCpe05HmbZoS+Imc7E/kmL/C7ADvPMj4J6M3kym9f
sV6woJAMSWiHAQPmJyBhSjKwZmZXG8/haaIRihULLOowU4hqB59gFxlG+wAai05r
+N+kDvejOKqnk+gFT2Beh5hq05AbtnlTlQ22zDTSKnpOB3+Eg/cSBz0+9UgZRiFD
FRQDsV6+tza1dV4pwPXG8XWt6tU0X2WAgvcc2uHV3s9VrM76PMpUcN1x6O8ObJg5
Uir3crWwDRG+YYlJjwWCdwj3keXw10Lfh6tWcKOsUOkPEC8BN9GtRLjAiMQO5/sl
LHDRlfYbIufwFD/F5/8fqEzJ7I5I6+/Q/ehtxlNS6Y4Zu7jFkKyOf4awJwbkYHGf
Kz3euGvYbmeAa/BGa2BpPXIFqzYiRm98/MuHNr6Cf8oQ0Q4Yk98c730QZtvbfLtG
sqCLe8Xn4ByukCvOSJroKpu4BLOBOKIKr8LoYp7n+HcgkOdeV0EbecX6YgGvth3A
MJazC4/B10WdZiew+iz+QeGz5QhZmt2EHM7CLI+pEaP4XOC4lR9YGBYiaQaOfb+g
lo9ecABk4ZYZeiOj/Piwr6pAvZyWkQ84P7qHv9BpViMIOYHxRxpZv9Vyl52ixL4y
2UbOJ/awI63DpZSZDsbWMIOiz0b5W89yS+ClPzGILG+IAToa9KpKx2p4yAn2Bl3Y
k4i4NgMYqCk8OQ2jU5/Ss+H10YfdMqkYt/TgLKl445hoz0y3f1jEPCjFbkX37Kag
/Ml8KcBbgLMAU9eNUw3UTjpZh3Crl1gcHyThd9G4uN+LD+r4iV+GHuSxJli85eKx
xXAdBEM1/+IPDlob8jjlpgBh5uP33xVLKsPUCdVPL9ZU4Oiotgew+RvexYaTnK+k
YmaR46VhOQHSJ1+3SoeIB7DKDsFePs0E7dLdc2SuwE9z8Aa47QfwZ/X8IK9wK/Wi
OltZqj5oMCGifm6VMuvU+MrsA5gq5qotObVZKhsWqKfPUC2Y/WvWk9w0NlIVLo4c
FvZiBS+Mn21F45N4ZV4hSJD5OaFhgB3URzsWYfJRZ2V/udPWBV6dIIvgG0WLUL4N
iP7JShO/+rC/Ir/OOw4yLKkWv/5uD0rjx2mDFMkXJe7kMZNOy+QXV9zhowEu6oHw
Muv1M13Js3TH6JvVipYAT7nzGK8nA6JrDR41VYOJNVED88re5QEoBmW8X413hO/F
+fQBVY42IqQlEapMtOK9v7Wrxwb4tFimlu9hDfVVRaK7cYkAF9LYsZeZrNj43V00
w8E+papu1k0hm0vFCCQU0GiyK4uxGQhW0ZLRzFF/M3DOZHHiiip3m1yzfV3GIlWy
MOmBZQ+VaIgyWc2+wIRJzUYbNAVvXsBiVUnlKsByAMb+3XmpzHONxYqwpF1j+Crf
R7G5GzRmH0YMacbHO/lmKkBvjVDhVk81hovghYn5+vAc4xLhbdf9lkxCYmZWllaC
ZIzezEfowmmzE1tOE5P+l1MT093nXuKA1aTUJBte+3JMaFAfyDYRtF1eHndXUgxN
fota7+qx8hYjYdVOGs96yDsL2g44IqhSSpDQCZ++pbME2/67E2RvT9gUYTqIVRqU
1fWHkPabgln9YEJtgaPI/oom+t53x3UAnrRxCTuvNgsPkksg3uSlMmD0lYj/h06b
ZyDTRgXv4qVlp4Q44OWQ59Zq7Aev2RTlY7pFdi61rFgxcA8+lTlPZDr6JhTJQVTI
7Rk9/YHf2bksd87DkOSpLxrktnhxB+eyGl8ZWLTYaRk5LZPtIvOFTkuM9hInV4Ph
Dy434WRrkgWSGtNeWHrbnh/IOR+u2A0+bFZFdUc0lVzC6mT7vaTNHsojhMVgmzFc
9N21NiN+wwqu/u8M7L1U4uHisvdQNeLVLpFp8VLFk8/Bm9q+m8Rc/pRvoInIRFBq
nJCcUzVUo9c2ybA9UPar9rWoCpyZ+iAjrJ5qHstumCQnBYnRpZkmyT6/yEVkX7V0
3bzYYoHMM0ZTcCpkgRxFpehmCQHVkXOLQy6QGLWI8mp3mvuvtXAwLgsw1JJ3uutZ
C3uPHvlN2RZvtA369oahXQsItV8WxNvAatUTqJeH+wb2Xy6FtCSNmC0HpzLJ/v1U
Q7kS1tVAeFfSTuwUyFbnRXjBih4hcJSA///81Bz1Z38ziiI/Ais4peiSe3GC6qiS
oO+OPGgVO80kYAMlkvUP08o2+7hOXCA3mKcOB0mVZEc/7kP8kdHYchGZZBG29yBE
ifd3htbpGRYegRv/OdREuCOx+vdNix3QAuhcKskS2bYEOaKJT1huWRkxTdV6bL/A
mHbVkj+wFCSU1QAl84IDS1egGsFEZEOCoVOokhFMqi43YkkEBEiLPVJKY6KnHiFJ
CLNnfJ4vg1pa/ijwzj/s4853+gbO5zFwyslm8k+sJMyUJDZpF1cQMj554WY3nhfQ
RhqV1lIYMRG50iNt1rJw02qqfGDGQpAfxHWfIo6+rkTROqRP6/y6Xd1hKM0Xla5F
x3NbxB9OnN8y6TAkO2KS/UxdCj08k3ZzMAaWkum+p+aqNVwxoJqPCYVCmPY9GGYJ
OM4p3SuIV8gXFuIVExaGzRSkxfpt6ENGFWAjSjhLKDipaAN0zXl5ucnnUDLLtSFs
5B0LJIw2rTpryAKMHUnmFed5S8aDGbaF/V/f/VMej0MgXGsdrFlogd/iZK5mB3eW
HiSyrwV5BkR0XV47Qa6WzcOKWFXlpfhFK29evlqtHIQwjQCncZdgXt8uMwvwaaPc
0DQ9VZZBBDBOtSd4eK6reJuYRdw1WZKFFSnoCUUJCD1uWbVRMxk3DSBdOBe7fxIY
4hQW4PcFEMU02XuVdr0/wh376tPdyHJXqDnY1fJiocuJdGHrSi7M9ce2qUiYSM9H
o8Zkmnofcm7xqP2OEx7Q4tG5tVqaEWaeZ5wccYmn6TYY4RWJXQLz0swAgFsob3qQ
+CRZkyxEe8A4H779VBWfoM6R5TNZL3ucnrt5WNI0M8oqb5olwX/a4kUg0lucyU+d
R2cs3AwAQexNLnFSmwHXLCm6uCWxXv8VVFTQBHgGropvI7w7AiSMV6eFpvBuymhH
1NVbVQ7Vqpu0VqgUwl4RsNRCRF58PT/69GfsNR3XivEHeapA4V68xh4cjXaH4q1a
Z3G5EwExG6B+Smmg/sdze2EoDj5OZRi8NVBVX7YgVU+QO6Ll7z/fNdydxp4cFSG1
p70LzPU175SQmpNDDz7LEIbum6Ak5hi+/pmfBESgIUxgvVI7KumGGMrxvMkrw5ND
/h9WK35MnSJDxfINai95NLNn9r7uldXRrGtNhM+7GNBSGS9TS8HOjZ8RjmEq008k
ztQDZ+UoqgTyX3fahSH33DkgvYwZRTY91GJmSyAf8vN+Uu9NSZHElJGA19f2CWEG
+Z8MX3uQUBb5EUSqD369dzt0fDnB5+C2EykCeHy4Va6eDaEOy/Kr3zmWmF43yoMH
URyEz4niaA0aXPc0HQTB1da0d771GLMiJLtloxPAPu9NAD4XJqu0BPIMOJKZ/Urk
bR9E3HkRU1AtYawMWKdKGKjZwiuFDD7NLvEDkyPhKqhM3V9PLBsttkuaQmRdO0C5
bixs/Dr6VIq4pALuAXe/RZNtB76yWi+F/cTjj9XcsSy0TB/giLdc9/wZX4oWZpCO
XbmyYNC5JMWtvZ0rvFcYVXDL048oyHphXETGQcsU3Zq1CDh1Ppu3+M2wGL7hLHze
9+nC3/QMiMWz+aBAjCJCj7UsYo7o2eOpZkhrO+xA69rgG7PXt53x9sAgDVzFRXB+
Bow6U384sPRz5knn0H9X/SF//o/CmfEhCg4HpxGGzVwujwXmOjIB0idufJhNASLd
tZCAhM49jIvKDH61ldunVNJ+7ztXShVDsHFi5OEj1rFqqVXiz81h3g7gWJFjle/D
s94+UotPfXujFQFAzS5k94JRrckd9uFzg9GVkfxl2YHpDtkOZUjsAhKsZlWyHj10
rg0ahbBlVKPliVcRmI1VEvbEXfQApM9CqCbENrAGLBoXn+palGLpXDgSMw5pIrxR
zxQsuMtgZm1YIo0bKToYUZlwFWx4d+ry7lqUZwu4EmD1eMzaMd5z8FINSyEcwkTl
r6HCf9HgAQ9ahP7PmmcjT0ZOsvum4HEZliTBvl8EE/hr/ZepszLk/v/DbBMsdzBS
OlxEdJLXIDZWiwesArrBw9s2mMn6COCpk3xRaLewqWTvZ7c1xZnLulzAB27wmk6+
UTLCfj73tR4la+5iY+YCwiBAT+zhC+AtZB0lKarTZYwcv9IBllY7xHE3boiENzi/
5ue3ZjVAN8pvqB7PfwTqMNo+JGuF9+ocdHjfAK50/T7pMO9YIguBmCDcq93ndfGz
TBkC3IJ7XQxZ3JCiHKLd4gRHFCOP+FQBQt2+eUSfYCQh28H0bjYMEl9eYPU//pI/
DpmOvvw58+JtSOmI0JFrb+MtaY/WR9iTFZ4bftMUNI7kpuBFcqitXNg9NH7wy0e7
Yd3dvi589bRmpq7AywZInt3tK3wUcUW9reVmCVh51MzmU88RvPQzqQB6tCMdPvQ5
2hAfc2zu4j1M1OXEdLOdOrXRyZWD46F+v+mrvaVYO1wzWnRHRVs7RFD+kqPdlcCj
FtTbF+kCkvpt+kG+HMEj73oxn/ecRzaE7XrWx0cW2U+imsCUSEYE/UMEnARPE2gY
PfkpvOgCN2OK5b7Qm9ELbS9vsSP5bXkC5rOHT2TeZGho5EysYSWbqyU+hl3F9kNV
QGV/kMdcTH1AKZp7RaDdOtNz8dqOg8PBVqM95uVIxHLeYNGBk6kG2geqb/9tdhsF
j7aSeQuKlyA31dMWEmml4au18lMUttP75MwJb2iOyOGr2FLc1XD2i5A1VlUF+mke
L/ldmM2IWrGMkI/YfN5pklwgY4yWlz6bzKuYxuevmWe3FfaJTeEAevApav9U90ou
Z6yWjPwFOj8vcV6vvk7/6BhuciWuQL7PD6CMeUlxgOnIWiuRj0v3AsmMvwHgXVx+
g1MPSW02ip56USEK5T029RQEVTEP51ugSETE4X5HT1xkuHbrbswQWGaizI16OuXp
LcQuvp3A+YaULLBtFuq6XPy5oVxDq4ay6g/+whilG1+ELqru8SeEZXfzoBMGyPS+
XCqZwdzf2jkWYjVSYOyqMENNYmTLpGseDNqQROkZcWjlKvq3m3ItYO8c6cqGF/jY
VYsrxsrnQM2C99d9dLsNfy8GKDcihGpM0sMqto49HxgHtbixryIMEofK9FHBmH3U
KN2C3XyO56ZchObvyMPf7tcN6xl+FynOasoqYXxUvVvco73KMOMNGkXaHXYOaGE1
eLxwO/nSyfW9wzBD4IHilykYezx4i+2tUtpEcoJN4nsMN6Y/udXOlua9g2/LeX25
vOxZ0eb+lCu1NZ+ha/noKWRk3oGkqqVOfJ6CWQwR5oUN2TXHaJcRkDlq0WN1nY3V
WJjrYVzGO0WTi6Z2W2G9dyO/8bMl+1+KVNUhpiCM4rrHVbZrbIPvBqcJ414pnLII
PTBkYXwjI0RErQVqr0wVheC5ONYiJtEYZ25PvupeEB/bnmGqhls08JGXvHVnlYoq
aY57Z6E4RHLN7878Qq/LcRivmPZQXpgyJIgz2iYI2uWwzlMdkOo++7Xgcw1XWe5n
Q2PjthIQOT6jl/a83TnmchkYve8PYPrVYBZLlITv/QidKg5HGuf2LUXMlnl4+Txt
2FGw91DgEpOBkpK3zUBEETuU4INQ8vauzay9TxT6beH9yEoC57DD2KNJoDPEwHmQ
lHdXlOIGabUH3q9+3KHOgcSxyUzxqTfWxuP55A7EkGyH9DXzeYieKmJx12+bDMOE
C1BThiHjGZUectB62M05zHh7l/mCLL36y4F3u1U0YdehsTakrPFikOUUyJSQiVft
oG4ThnRpQ333ZFph5uUfhcjx//SON2NsmpKOoccQ2IbptQTUN2lNr49Tdm15qefF
woeKfJr2qoMMIeLzCjwFdfmQqSa2GdMh5iN9fRAzC0iBIPXKB8qcKOpXaKCCnBnX
j+xgX18a8p6mfatAB6p3unxJLMbhhX6f7NbHqxEZbjPWy8sP93DdZYvJWMsKYWvi
hVVQhnSlIl27on4zuGQYTrT50uVJqXdCvZ8DxYPH68mPE2zWs/SNSksi2E0H2Z4S
KGow8JxCgJ+s351NEp63XLe1YB3iQw5FBKuQ/4WEP8wj0q4VX0KDgaW7jNHHtGIB
KLEzEjllMoepwxq9muO6BknuvYv5wFx0SY7UmpK55M75veo7qzj4HgffEr0LgYWu
E9W8CdniK1VNUyvZmui+LHqbiCEcG624M3gMSQV/soRwh9ms5Bb/lQjIzl/n1+av
4e6hCFW13bsAhMp868jc9qMbNsw6UHAHo5Ndi9iPYILIEdbxv7t3n/F/MRwFKVrF
aauPexU6OOfLbS0MobODlIZ5XBNvL4ahl6HcGClYzowJkRjxpJq4V58/upKhPVcn
JV1etadj7oQWhxgiNXiXaYBd3vD1fY5fSH39lqGQHiwZt9/lnJtXPetxtVMQoPnB
IEFBsdKo5SElZfAR8SrS8wKZZkzvvksv9n5iXMQyIpgC4mistVYVwbhGVVn8ctPE
FABIfzXTnsY6KrIqq+woV1Xci2uAoPeJRIhX0mErJZhJSpQpI2Seqe0cpbmuW51U
WECAB/FtLRs0GeZT+qEl36DkEj/qHyepgZf1bfOqsCa7hL8YRoyM3QEOH6+xgmUA
Rw9OucMVSzzCQ+UoqFipkOHt3NSKTTeepZbqg54+5vSPkPx1FtLwB+yEqBp18l85
N89G/HPwgZXI/KVJjzBKxTchwBb6b5VHQLuBeSeQYwb0BqLW4fSug1m0n2tCaGHU
/EO34Q/WDxTNy4X1jwa0WfQLuEZNnUZCtBCHk3B8YPe6oQsR/RXO+umOBqWsIkHm
ZWyQA9WUQlIa4w8vgCWpMYdU+trr1jNz/ZNgHozpUcMXqkwWyWYjpOPI/PImww8K
ZmcSYatIgFIFoYBIfDv4EaF+fAxywTWx0R5R8Q460zGZfa5hDmi2/F6grGC56BsL
cjbIoFXuZtadeqT4NzPlNkokpcid23rDtzIu7rZbZktMxevNZ6lImG640YA2QElG
HGsknhOtvRg7aIZhF571FkCXrZ7oEMt6Xzw0cQLN7wT9vSUlOxj/UqJXudLqSY+V
s7bRcc7iPFcXwy1H20oycOZLShOMmhTIXGKIdOs4h4T/AnQTrh2BIUb+aafEjm1r
vW5AVWw2zxGtnSfweg1M6BSPGbhgOnpCErCmtDPLw2QA2M4sKaEamTGjKG71brIZ
vY/GWJLbDDcXHfAQd6ciItBLbv8R81C/VeUYfNSZDoPEHJOJ+1JnoaJbdUweOlXw
T0nrapKfoTngDOSmz7NHS8VG0OSt/9AoQNwfivSsfLY7/3ZizQvkpFQMj37tY3Xy
mvYc9rnsqzpI6sMcT0xtZMm+VWYHL6nC6w34C+6YA5fKYpQQ6DgoTPBuzjIsEniY
P/h0jS/AH+G/vfn0noQALqiYJW6EGDxCzLiCuYICM/UwtkCYawMl0qzFugEYqIPs
nOaTUzYmWJyGZDqh6k/psoq9BK9ZZTTX61REivOSlGpBHsLd5MDbYHOy1TJjuK/d
B9U8Qr/RFQXnysz0jyOuBfClk4C73p04wryKvxmO/9OfLuvxMxr26hN1yhb23EDl
lbPm3GUvp+F7OV475gd2KfLhZdO01/wZW4hTKokqhJ435Y8R7RzTXa6dQ6UfC4UI
ER9YNyg19q2k5mMGW7DGbGbeaGYp10nMwPLpXErpS5SSlWtJjiy42ACvWFCfXpqM
78vuqOGuBqxeRX+YT5QTao8alGLKwbukdLkTqHkeA+Dik0oxRC5t94lL8EetG2TK
T0JEOiEmYdz1f4Unk5Tvhjhs5xIPtHPbj5J+aafcRkyTnTiiXamzp20jadIxeoNo
kkMx+zetzA4sL11l3J6Jhs5+2s+MICaGwPpTp0zyXUhigLwJ9xhCn1g40xI0LxNU
m5ZA1dj/hYEUfjpQ4NLAnOBLLNT2sqJzZj7Ye39pWj+0BWF8ikTii/CG6ntTzUW/
mV++0bkmiQZpEhYN5f74as/r05x3u6r0VNJl7iXC14+UgAqtCtS38rJtPsa6wEAF
KofZK3Qqvg2ZoXg5FdWXuNuk90ojCvAAFOvUYLc48S43HiZPFLes5CHK2Av654yO
sk2AZ6NCPORGaaOc48zXy5bWYR55YQJj+y08Wq1aM0uyp1lN3LmkTFyNmUFAYgbJ
/MHc6akcQWMCO7b+5l4TVtAGzhZGbY9WuyGQdvpaCrHfUZ/iVaY2DXN1cjxWz58L
GPfUDmYRmbYrBzn9KhL9VhPWQ43/SCDC6PlR4tg3iz2MosGyhSdl1c3XoCzTidBd
joQNgeqWgGw0mNjHUARHoDz4crb7s8QYUtWgS0HGl8VnisdAo03E2kEBWRqIYT5L
onRPaiHJL+9XGz3LluPMAN01l23BsasiCo3pYvy1jtINoNR8U927cwFyL6HtH9ho
clk+3JhDit9UVWYojOQhpKGgtFmZTnsr9eJQzeRhJNlkZFhQ6wrgnrDIFy+LfZDi
lmMjGAAm4kXgz9M8CtzvccI5wSDhQdjm6wVVXKIcLk+Oa6LktS1Bpw+Wb5PnkKIH
Z6eN96P44lD0FmTCHJ6CmoJtVvzNYQZ5VG/g6/vM1/cFdVxsAl2+NfgW2Yj+o1yj
Wqtw+ahMNFax3TvSip6JmBcgcXPqCCkLR8P8Gb65VRBgfDU2vgg9wLmrn8XgAVxr
LkBFZM0IXjR3Fvxg8OF8rIKL502XzMa5u7Zj5RdQL+QBBnmpWhVTvdN3WUjyilzB
qpaCK5ConC4ke+iCRUm8JvqqYCchog3gfPYfjOiRMb9VEuSJZ+Z4tSnLrwYuI8XM
nI7xrntcx6U4LRJKszVQB3oIL3sPCW592H8gQEKFvMQ44QoZHQOEvAH4rOQwg/5d
vJAvhQxyuyO8Aos2g3S8+oDovPjzf7DW8bECiSdDAnTAQbnJHPqwWF6AaKDyI8fw
BzvAOFMpksb+KnROND+wR6ubksOYFplGpmcufJYUNFb+4FfAJC2ewSV81fqHPIap
HHLbJOLoOZ9JJRMbmbHdCgnqV4F/wCVIAtTKMbGetZb7BMOKF11zKdqzy6AQowME
/85JPRck1SHk5pf4njIH9rrtQxvNqX3yac0KDePbuvWUaRnqfSsN38RWfqpiKWo6
9KnmHJSkGN3lWCSsp888Gr7Qyc/iNK7llbPdWCalMqefzRPnEt2NbaLyh3zx4Qns
GJ09fllf8QJY8hChJAcKSRDA57FpYG2BBq0Tsjv8R62Lmky+akJtCMVa+b+gv1j6
3q/6PObR4UgSU+Rl+rdVsig8RhZUsq383DPLSPoqG61SGCMWFzS8tegjKFHxreQX
7TMgRtMnuXfcIB8diKp5I4ck4W/fB3u3O0PkhAdmqfWXPl/m/1rPIPJk57+E47jC
/xqcKsA0U6EArQM0dq2oGzPrf0R0XvYpIg4sEI7A2Xs1iR+UVzF6Xkds/JjVrP1C
4/JK4go6OQFGsetnBwLuPNR2VbBpSZmIGZAyxZFZre6ap9SMI41hW3i67Auetlvy
Ml5/Dr4wmBN4/cqvbig3hl8iPq+rXCiUvF+mWRpwNA9OZQh/sYw2A0wUFYhi6CQa
DuiHd4Jt84MuRvhBcLI5fPXxVUiBdJVhd9DdgfhZLj0POsI8z8j0Ts62anV+Ng+g
NehJOy5uUEEo+7CS8bB3Vre5CqSJDC+LN75NYaGLhcpe/wbZNkYkOYI0zThs1SSR
4qvFKDqNB8zn9f443jSzPJFeTxoahVLrfzxbdjy2GWLsDKIihOY7Ky6D0Tb7nK3y
9FfCvT6DaCGPUBTSZB9v2oFycImRKsjJgczqPsbQ6TgKxhL3ZKXhJFTkMP0Xs/oY
b03Ht7Nrqm/nWlw2IUl+r/IYjvd8DN/q5eESI5aMTHrqxMdckErlyqI8sbWWqmV7
CHgMEx4eGnyzdwVm5iY+3l3DP4fLbbwxO672UFbM0QHzzGMiTy1MQr+lZInohoSX
yHzk/l3wa3hGIbS96L7tpJ5/6F/tmXgd/AgAebzXTwfT9E+IXKjSR08AJLMU4wI+
r8ebcbh6mxI/gp2v+gFP9MhZstBZ4Oro+PIz4yEu1ch/PqJo6EfYyH3VPvghoc0j
EqH4saymtR13hViGxeUy8NERMMzndNOi7Jdyrwu1RCsfW0a/BCP33xTH8n4dpl1L
BO9ZRBQ+HQc1JUIms4+E6ojv2f3qFZcglZyIrWFbar8O3LsPGkcVIPPyS/k7QBfI
iKJ25skB7mbci58hy/c5Ku1Pmkihj6cfMXA5YYeId8k53UoxmwwJZ2cflSIV8HyJ
yLR9aTsDpBzEzsYVuhx4xA==
`pragma protect end_protected
