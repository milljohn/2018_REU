// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
E9r/cpTnpDidxuuQItHjiNi/SseGbBkEFKpVofiKhTJe5g8+uaAlDqNdVaBqn0Ij547Hk6PUBTM0
Dx5muFOKb0w/1g0CPE7D6MMNvQ7gC10DmPKbBQNr4aCXPpvH5dGWXgMYZMjhru8pGwCtbxlY7ryb
BkTWMROzITwCWcszvyRJLc0ajT/YWuZVofszc31eiqRBYmMeUj6tSfjD0LUOz/bbGkb3yMtZSPki
+ToqwA6uqyb5Tuc1oOwxC07g2PJLFp5VkTj/uTAhRxJlYE8DjPxg38aw0k0auqKh5UP59jMbh7WG
Y5F3EyjHGi4uy0kjR2Cpya2N5RktpSaLjuImYw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
RKwUq4muIusBkPSQkGWh2IVFckXf9HrJesPqgeeNrhSQO2HxR21x8zmDHUsIHTxbV8OSAjJ2PHT0
4BidekYDcPURvktXKYyBm419rr0n8oYYaoxL9P9xY2mDXsn3Wr3nd5Hvy6cYUiwav2Hz17Yw2J6E
+h5Hj6GYWnAf7gVlqUCF+VgEGOUWQ0RXVYuHXwzhkCqVRARF5cMhu6hm4WdVR6E+Ydmiw6fU4tMU
oXAOKIvdou0Ms5C4womkLnpuvUogpbBLXvlUb4AZwzCZHr50ac8gT+pjejLv4VjsJrmXvxCeof6+
d20op2TZG92MTzvRZKYX+dPXKbIGr3MU/PzQR6c7RwC0ktERN72W6M9sR7tqP4Vukd4CPGIX3w0f
OrWlPSh6SOe356nDOHOFFUzJPK2QRQJUC/N79/dGd+H6fpQ79+BDO6XSeB0X+V85FVzUjNtNiEHj
sUZTMuiL4qu6rA3XDUMrG1+Ef62G9JrbiGXaF1GKdL0cXjxBWNDfDMqnFgWdtSXva69TsTJMT2Gp
rKVSs/zBB+QnfNRktQ2RxDje6x5iF7QS8OKfZz7Yv04WHfQSZN8nvrazrFJLCFQIX6pyLVl0s80Z
eYZbGdsM7i0lgFA1apDySQF29Pb5WLM10fHIs8hynpcbD8h9F5yrb/KU6QuFXHBAGIbBB4GS1un6
jlWUfGKjns+NvYxvu2qCvOPZi/NBTv86YJxmli+nmB134Wm2qi/U/fpJY1nOb1ZkT4C84UcVPO+k
DpTwHq2Hg/+Orb/dvjKMeDtH/W5fBTAdWJ0i2d+1SikfRXpsyMXoLGNGOtj/w/LFKpLzEHYtRmCW
4DFLAoZcpK7s6r3H743185edJP6bBqSDSK3p3zrlbuCCuw4k+KKSFfT8ujaehedRLOx8ssd1Pea6
A5yAThakjfT6zP+5eXo0WHgKCg2H30+mT6UtJcN+50NxFEFGQaNYqmKCP0Xwx2GluzTHnFjhue8B
cpUgkXr86kjRr2dmFLfcAecyejVdDjzju9tRc6hFP2wKsFJip1HP+8hplUQreg2iUPjFCik3Lrgx
X5rvY6wBztrwqxWfWOL1AGtU3GfEpEpTlWyWFp882tiosRDe/xKJzosNuTcqoRxtR4meaX0hgkYm
sE4RdwhAFBM2+40iCxrF9WJENtYwajigx+GItUATR3/Mc3DdMZQl+XAGAyq8VwZWkj5lkw7LtTKe
nsXACrzvYgVTP7ZytNkWGeolLWzRi//5ZinuIwngnwcU4inY0IO/5evlKn9WY2ijk5924GcPCphM
BnR7buy2bbxGlyp/VeFosFpqsHE5bHKENkZ6eye2QaDk8wchptD6TL9JKVaaq2xwuMBKKMyfZANb
3iSeWGs1MSnmfdW2uD1Y3WIf6eTuPpaE7mk0Zmsl8rPGlKAWlp/LT3xNzcJ+jHIcfHIJXywWiYEt
g5zde9i//kgHs5h5bGCjxIjdgCWtJbWte72T4n6lS+OOWMjfJXKgnQXC8zsaR7bkFwfmgcjn5CtT
P59d1+tkJRjm9fkncXEx75H/pONMTbSPcvMDUeFymkQdiyup3Okqc50zdhQuM2cW/awK2wQUJ//k
/tZoK2QC98ResNmtYOu5vNzvMAZF7cn2V5AjXTKKz3MZzebxsT3DQlpioxIgS6eOkUh9iuNAj+IC
T0XoTn0i+ozN0JssXktD6YN8t+8VfeRRNGWWLq0SD9Zwxwd1m81YbZObJdNkzK6byMr3CAy0Lhpx
A1+cGI6dUHgnW8n5rPnJgKNh9VrpByVt9k+mv7L0FQHtIdjpe7cXFRdH6lLlPX258PZWn1KYq4VQ
AVcGZdk9V5/k465tJAqB6hUCwQ3aEljfC6YpCH6VIh41i1rKhvmxInErfMSgJPcrSOvpohI+DAt6
zXVC0qluwjtAoY+C9qirJ+N4+BP1IC25nuV8pQROFdJTgHq6OVni2qQvGHJjr5zD9wV/wjPHk4eF
D4/8SrBgi6BEBOnQ5+DsOIldZZmUkEDQQMm9KBVvRnMJYCcbjRbJ0CMhJ9dV73dB+NzsIelZVu1y
qeCZT7i8ZInqMg+MSSts9qOLu/Adt19Pn+ZM7334GAPHO9/O5vyrU/5/BzcDieBWlx7JBW8LUyK9
hTqqpfOVvO8jftzS4GVVnL4G1glvFUxtLgLeb2z9N0/9iGMgbKM6ujZ3beF4wZ1Qg61joCvGK5yk
J9hsoaMLjU5kucDPYEDAh6gziQe0xfkuKNi2mHyr4shrmZkiOuUNuXL6+FgeG9u1euQ9rr+8UY1T
Ho/+yqecR0cQ04+qrZ4+zaOPaD6Bou3Ar60/iH3t/hpn/uc+sPr9iWsCuQMYWlb5gQFpC3dO+Xc9
2DOQMCO3GF9qmYPgDfR3jIxbBz+6Vge6y9h+glouDCXqKfcert0Dmiw3b3yGDAF8y00Jgdvvw/2L
A9DDJu9GoI0yfhqPcjeVP1hnegfFMqIEYbH3LXsEf7JfFEI7cDaVEUXHR3NDRSU8dFwXZoyfJEMJ
bQA00fCZjlnpJAg4I90CsSW1nOC8XPfjL1uSU0GyAHut9NAmnHtYExp2FG/ePWtb7SQTtiSfMpwI
r/y1jhLoQAkZ8Y6CqK3DVpMQjGIetbhh34MruMy9oos9rBd0eZt0q5cIORdMfHJjz0IAGMCUiMU7
bR3+msh5qTQlDgH4Rfivv5shAeO7PxBCdjk9CMDSR/nMwlt7UIlxIvDYmYw/olnY4MaM4jKT5DaW
Yh2H2ey8ZZ3W/sqbK6wtEUkR7N1pcLn4KUGN5CHnNu063+HTTtmiONqse2ZFDVdyvFllDfSBJ6Zw
PV0G1+kAnoT0s1wYWoh9yCisVkyCwR9uievNCaof1rfKWrIMReDilCkrCYd6gLdNRPNeWg5XM+5p
jgL0aq2z2KWKZ1rEVq6e/pyu+nppTItq4L1TYBKX5iLT/9HMGt21NGJg4DZW9DwHBV0RSc3VnaHU
NFoGdWOoqvdT+xf1EYJGedasugRgJr7/v6i3NXCLZ31XcATUo2cv8seud6m4j2PLVSBUMsqxqYa3
L+uFp8eoz8sK/82Q1ZrcIr+ysRZHvF73gcTJ8iXt+MtE6ffd10kbMeiT1tmkWVDnK30AdTMrykgo
61T31bX0qDTh6K+bSpZboJx/Q+7mQhwkXKO8mTlsiTEWngNRWtGCOHpLcUMFCf19M8zWGVKYuZSQ
zxxw5Nh+4ebK34VwiC2hYoFnKOfrYvB3VMqB6m86ViedYjLdXxkgb6F+OWlGzq3jfuLpj50qUwf1
6M1cWPXYoPGjfKd5JwqQ3uGiIh/srVpYx3xHmkaX1DIByhpC9YxA6euJ56KIxDHX+l6ErdkYBr+F
7XZfpgeDdAn9+xRzv92gu0f5iIxDlTppFVlD+uFjNx7UVS01Il8JVw3BhTkqHZrlN+RTk8rfrf7C
8/bVELJeclrGV9pv/zr7T/EueOxorFgV+7R3uQiwrgmTOMG8mOQg3TtAUWfxQQF31KArp55G0aBO
h9FHEoqtKqpwr6mwH099DnEcanZx+LzHQiiRfsNYbWHpTDDC0OtDw1jCKzgllV00xuzfj4OVsGpv
AEcNHzbRFvEwYz+vDR4QqKYny0PgRLEv29ndDvtYHySI8C/VBjJKwkbxuvGF62BX7mFbAfYRy8fI
7Omzj4EBauQL+1Arh+5UXRNW1GqEVZL0aDWJ1k2DyDCZF0kn8ZpmCo6joHmnYKth2sup5fhL/342
aiTABYSGb1KIE9yVUZNwrIAp1iuDRiETM96RIXFNNJJhvpgK57PWE5dm30I9Q8l7F8APK8JleZOD
d83ee8AHSF8AAt1RfSVJDI76/gBnXykDiHdGozrokDq3Crela8N85pK1ieY8stPxAvU1anla1Qcu
9qM0y1taL5hApuYXzCVU21UKdwKA5tKHP9vxzAzejHI+3M6v6cZOxJSBFAo4TQNk//71bVVMIv2B
a02Il3xjDBwDaM662m70yu5Ag99BzpmZF0Xu3CUbuqSqHwyqCQwQ68ZXgQMUaWtiaHcBOWxTsnuh
ak2Y6V43YG4z5xXswuwthgIRIKqM7SdbUfV8j2EjBThI4ZioKAolai/USVOsQmOt50QP75qGPZgv
1CNFpOsIuQFZpn2mLny4Zio6MTFUGytWQLZM609BsiNemKxLTOLyinYUQo76GHOvdo7/cbOp5adt
bNswSwWxG2/jSo25cD1On2eqTQ8VxDStapAgFkEDODx3IT4HKKMTxKGiPkUrqFvZ+FtNi4nlEGv3
m28eUd4/qDUIdAiI+OhXjygoczOr9OphQ4hhMtdxgNlkvHmtZlmSP+DYBLp0K3yYIeppdcgUji+c
DuTeV5LaV0OPiRyExQU/2picgvbXfsnS2mjMNfRer4pE8uaVPClRYZgiIVDApc2dPni/x9ZRmv78
8NTY6A8Mn6qdQDiWgE9ESWnKT+PgFLP4+2Xl9YZzmLDQcHgD1UQN8JFiOCiSSlFkZJc2G5EccnbA
kTVpMbMVRa43bDYroEMF2YQEICw4sE+swwazO04giA/TygMU9ovy4rfb/muta3RSIC9tKdgiOt33
OnHpgHjYLmb+7x7QywsBBOQNVYOz8T7687TntVil+jyx5rX8bD5+ixhOYu8yDHTXqeTswNXPLedw
voi+iGOh4XHDs/P1lZP4FAk7E8d4Z/OXgWbS9YeB3ukaHpolCO3bAQWitQ1rVl4J/3VmInn25Jh5
sZ7TdEViF25iRcV5ORv+ukDUX6aPZr/PBdUoYOUfqO2cK83bkDZJ2FEfK3pjS6pW0zAdSbPVHh40
KZ6GlupYSizlSn5KFVOmk89ElVBn/fO3awnQEq1APVAvG5PQxmk2S9lWBShzmeTJDFbt3P89qE4+
0Ls40LfftTkhBEEI6aBqfrE0Q1G5hTVXS5kC8x6iZpOVJl04D64uZZ6qsx7kCZSOQJhHHi5u/dln
mo2PXz1raRithdcpw7jCliAGiO9C2qXoGZb7iSEwZniPGRYWH/qwMnII6kn+flfnKatQYpgpPgxZ
temFx+BluNCaPXvMBKsTHLQ8PPij0q8eHYzFBCkhwmApPKeYctWv5vD9oEGQXhx4z9ya+Sj+0uMd
lXkMzjqSi5npdCk3wc/bcBLybuK1dnPge6/yg3ikABrvpcA0/5uplbNCTCMi5CAOBC7RWj5Z8Ua1
IfnuGHWMlx9IwttpufFpsHHdcILpQavcDjYyZrrhe3KGR7OSLq/vuAj9R201gOd8xLRBngKNpqyd
nOr6JzrHI/a9l0NiVCSsUXoJV20bNs+hzXKko13OBxHVeAJDVjQZ2LIeuYp1qf48ByJbQPcLZQ4z
zuOQF12bqPIOqsYRuhrRCFIZtiIUfPamBgCaau6KfWLOwmSYVRA99sOu7/9FrDeliWSbHWbxsPJL
4/yQXagtdaP4K/SA3Ak+aFKzv60xI7Zh918j3I2bunfSB7L45ZzavzlIAzJ6zM9Voe8yUsiucOdO
VNXQC10whPr1OaADALyN8yD0wvV47zunEpW5E+YUKh3ks2i9wVASWZ37yDW2gUh0aBSbpXiMKSKL
K7fDqXGymXTvGA0QgQZLWj70Rebc+8UkKdi03AVbkIunKMSXj2YV1SEUw5lbKatQkRd8Eclposd9
df+nb4gWl2xHQJ1wbPbJmZN+yhoI1cQqeBFChzEujjNwKLn4wv5GrnFnCvDDC8Ds7DK3gTHFN7zj
8HaIIKp1YeeITU01LDl/ojXBSxcxjeqqGJl2D82O3x7etmhx232CoRlGfhAysRUDkSYxbb09EaLN
azwb/1f4ezkFRYos3CYDt5KAPrU3ElZcMHGLHrWAcvNI1XHZWqUDAfgCAP1XDV4FxC92U0yLZXDA
VjRfTiaXsMCowgceY9hNmsSJ/fuGCsxrnOh/RqCILIbTgiqXLS+QuCZyRHAl62lIUwQoLc89HmgW
KwhWau0Ym1qLRWUaAtz8dS8o1opPbo6/MtKMu/4Ol27GyTAmOM1YNsn8/yyqFGTjAIz32hMS44YF
lv7+x/WpVNXDMu3ZZkc31eT8EeXXl9h7noJUTLWZpOQp9F0fR/nDiSkMykQ2FlGwxezOz+S6FlE1
Tr4+6Rg013alUaRagLdMQWyXAdA05iZWkSyqHC0XR5/zo/of3jaAU/1jr5oLubDY47qqshIZcjoB
XQuMliKCHlpFlWqb4fd1EOPBgcBQxJdO/cEOZcgdo+6qcvuOhfuqpB7ywUehk7fMvfsASHPyHQfD
SsUjG6kiDl5CmpkwXDrvkxqW2PlwmWsKmeP/eolAjHpIUmxe13cEbHBCYI27+GzJX6c0VUGyw7+C
fMoG7gIKacjCn7Fi9X+bZ0B6ZUaPGQzgqSKq9tSF/vAzU81rO/mSpq/PLhwxzxcAa3aXRmT8ftqu
qyeNEZWrco5j+oIvNIUQ2E1DVn5TdECl5aByr5lXJGaNYHEjNkhNZwuh3z3nz4obBhXPJyTJfJjn
zriapACtntE7XSrzrtDFy8NK0dYnIbnKecqzCZYH6zf3uX2eV+BcLLoWRkUgFnVY/WPyuhWyb7O9
9WgZteKelfp9ZeLQJ4YmgvFeoH8ofC0mMi0ij+RMzM4fO61VZ/ylfGVPcdFvNtk3TdF+3WFoijWO
FUYGwR8ozc0sJ5pCMQ1nihjlatjmWIsY1Lc3zSAsuQyPS6JUyGFgvuY+RmmPV0vb9ySyo8q/VrHc
/8pjG2LFCwQqQ76/gjPQ2MN2i5yKOcJ1oQFw+fHc3hqKwAJFXML9eDNL5rnXgTbpTdVj7KvanizR
n7GBgBe1/S6VXUm/mrFCRf6Avc/vlSxy4Sihnt3tELPTm6g4uQZjmmKnWn/KLh7jiM0flgSQuyy6
KrYc42wGM2234FoAZz7h3mpk6J1LadHdct8lgLk24izRPQRuf+CMwFQt5EJhwvMspu7Tb6c0ZzOX
Tc2GUkooNVE+6FA92nuPBbRLvCUq6r9dn6K/Yd8jBp+NnJMIdEwRzbZU9EsyKjL381jd+PoJIlu4
ejHX01W6OMDRhbjQPZpv5asHSM+8Tx84HoqIsHdbVNqUz+R1q3cTOpjT4sRAvWHnGRws0rTwkbNR
nWvnBul2PoY4BfpKisDkaeIo/x7h2Xxh8AMu9cz3kNvEE+ppeZwmsxsCtEzHDfzmDd7YuPvHMdgS
bcOt1rayyHsTTTCG6Q62dfrO3ecEugp5xxZ+Lbk8Dqz1s3WDOi2BUbIqHX4xW74u1NW2oVEYbHPf
EefvJgc/lV0PgtQy60Omxy3IaTZ4bnUjvGd72vY3yRS/wnoOWCkpPQlj1EDs3uMj9B6tV3zHZEAo
yO5+XklBtQcUbrAEg4eYKYPSR2BEtqatlbJy245Vs0nRezrZ24xDp4109cQVwUGBJQ5++w/lmI7e
BaSQnJOY3/Pj7yHJMF++ElIDZuKoaaTj9F4LB2AP/LMZJ5XclrLu0eugrsSqoxyfNQMKhJ8nrzek
o1o7tbUPyxnK5mCjmOT4v9HK3qx+FyQfxdCsMJ5S0x9iAyOa0fSYUHLlCzXBvHF7MeQnqhA9nAzo
xRIsox7OI7HX8R6+vD2NvLaycZmCKTGrPVklWFz+oBFo3VfK/sGUFgKVLMU04NlC/unl2ZSebp37
HHc4nAmua18CBCniPn8ubajY0wXf3VMy9FJkfYbFbWGSYlBmxxMiq0cncDf7Yeuw8Q66PC/21r9r
/AEZ1jwmTYYhyr9v9E51X+ueSnYrcvb8zX7D/aF6RNil9jy6Mw7dH89ZgMdd/kyC+ZxAplsjOOwx
7DxDIJQie9Dg8YxLshIK5f7tqrmw1CZ8i6U51GLveJSE6mK1MS5xnWwAw65dQ4RIXXNrYN5dCaBS
To/NFzYv13QpJmkBbx1JGSRB08fTzdaqkeKKvOJneNa0ne+QNvHCobufUHHs7pYXD9rN+vi9v8EB
HKL5mXxEpEOGIfvGLcTivrhpNqwZ7m8nMS4rB3BEyteshjZY0av93JM6IOlicvuIvaeEx49xB3XR
oUaYEhjOA/gzA0UwVKCwkC6AEP56BLR30EURB/OADOLXGnJ8b1JrQ5UlNzdtto0fG1O5RigdOZld
eQRGmDgJPN2pkcGWOrvLxSHNJuuQC1HwAqaJP13jC+by8d/89k+thq8YUfknQcYZw7styiRgZ21z
5qOjWb5iN8TZ5dqGanAU6T5+ETQj4XBuvOkrkKBz6Nd1ds6FlFoq91n8t02TJT+FsTPxatlRFtrm
3D+zDqeC7pycHtEWQBKXVlS5tsBA0Fp0UJKWzkwFNFsAQc34y8qYdEsAViRb3E/PDW9Nz/GF5Y2K
lkhHeXN4zzTIfoNz4wHtxBKCO1G6BRGssuENDxlJ4L3ZcipnLkSom+5PdqqQB0y1TzSRf+TjhuV4
q4IN4vq9/nEa+E6r+bqzaLAgiwbl5df9O7NZnMFmZwJLBLvYaeliN9jjnHGc3fjhF3woA3L8fM4p
1wvhCJuNt2pzhULdWYx+mNKqUQKl/T1VvroIMmsaAeMbSH+kveP74AbNq90pY25713Opff4LeOE4
9/MqK1HkUXpKp9jXRFI3rw+6igyCxeb9V/lB3sa1v3C7/8/oeFi3fqd+Tn0F0q893aPLKNFi6Qvm
bw/DsiUs72owTK+YbeaKpXMqmwTgee3CIXD1///fFUtZNeWPMByT3rPOBLk2uPlL6eSo4l9G6IUW
iFATIpT48pEPrJh4Qz8i1k2F0aQjNh3pPA7ziKnUy8iQ1IPSccP1Xz4NE4jh82dfTaJbElfEAPEU
+8eGdOrZwVjsEbDXg68W5yoOaJDne3uAXuAYYRG2ZHTqYjI419nPMc/puo5aqxGjuivmIq4+ENH7
Poa0nQ3d3tlZ4cfSUMlTsS0tXk6c1AJ2lJZ3zOwYUSmglOE3wmaYH/OI9JCa3xmLVj+bINcliK5S
UeQWISETscfc62IG0/RsYcHk/QBKxhzDXqopNa4GBk9EPO8qASQ7l8H8s3dP8mNn5ai98rPMJ7Cw
96al1PuHaP53oeZX5M3cChniqbd1voVF0DBBQD8aDquwyTBsyS/2CBy5ofC5vqpnis7vFO3JCQBK
YxLpGz2vXVQYNCAMrzqDzBba+boo9ZBPCHl+d3ZEKMX9IGpEqS/5A4ZJIWtDe8KCPeOtJH7vYh4q
yekm2tfS7ImcIo1n5EnE1soTIcR1TVzXVnuW5TOeLdqwuORz3+W1E2ia2vPvpN/ZxRoAQjds/xhX
JglsmlifoThNgzJGvH8U62l02gfAmtFgBx7Zt+m0AIvakEABAQ8xqz/GhMjZkqgZlRDcXrq848m2
PZstM6e4vdKdUQUPhXacX7Hyok5vV3OLRMrsmq/7wPAFAC3W6whuQ4qU86AkiUtcsv4hbzmqFu8F
SEZ18MElDsHFdTsBYm5lXb9lMOi60Hu2cNCxXsJ+HTjromBStQehMqT0OZUAq6CvuQdGDgrElOaj
BW60yDjEcIGhmofyjW19uPLxFqGHdNRCYVy6mSr9FTV9eLyJNc6N9LYF6ZCFimQEUV4Pjz3h3V8I
NWUceBHugPtbpATXYuGgdYaCOHHh0OvfuLYKZmLAfj093wMEChz/V8or+MShApR6AiT9/rBWL37z
HwbYjRTkyJHH5uJ9UUS69decwKagrdEgfJ7ZOmDx58puUYF5w15oq01RAtVVdSRRTZsvnfyApd5y
W/bUMssKqZLqD38jwH8LF/5rr5vVY4CObZYiAKoitD0BYxARlSVEJ+OUJQdH0t1rr5VysZf4rBFR
gE/ZOya+TUXV5Xe4Zef1vMTx/70jlRh+jNZUU9EFYCNfDn7Ta1wOgNytlkOwT5b+blt+Vjq0+uj2
XcjLgI9BLFQk70OccrrbaLOYpSBzAT9kX7xhwJSVZ9pmojCwmOFd5rDa/irkCLdhcI1lZ6FknOwA
/eHK5DjX0Dk49lW4EhucVEDSl3COyWvKcGf5LAd2sPVkJEWIIltcI4pVZTZWOtjNj+mgDsSY2uVp
2JAGgyfoPXNNelJZkNuSTStHhJS7p49gy7qzeiHIAWkpO4vcHrxyo5jtmjlu9dkFHrRkKQZTIM1g
94kis5rJtPocwVGF8T1q7SlORPdKB2qVWNNjXvcJLswxlDHJ79gNffQxqATP5zQp6z7BTW93D55e
3cVD6cIEeg4Z2lCV5v4EEaNhDp20bkVo1+UQcT3kJgGxPBUbfpEjIoVu+X8LJFkuj1KW+srSB0uD
G8Z6czX+XxKirDMsoWHjyQBAixBeELtJXMRAE8rmMPOsoFKmwF0e6/BHCUMY9ZsgJxrMELN0q3N3
fsDrr8Gwtk7BD6pnSaHeo1mQq0Zwu4PhVjTBeUblMXITMffD6+3buCzUQJb4ix+fE9zuIVVYSsNU
z+1WxE0BbmALgH2MSmtAje5DYNsOt8F8aooi0BvnbHW/H/xUb60HS+X70ze7lxMVNb5e6IBSi6vY
bB4I8okzz1QRCRuuGwf+RXldnWiyI61e/nKsuuG65gW+mpGTyOChZplQbFEfbqWtdhZHNSvqC3UL
Xbwhc6oCj4W8OIS4tDRtD7B7eACUfsdHgergFPrwEus1Nbd8YFBdq4rdOz4P3VIaxvkiBazskGh4
G7bmQqbPz4QRlQxg1zA8qqxz9VaCQgzqdXHP8OctD87FjtOpHcs40e+lqlk6maKLslKxQTsyNn7h
8WEpa+Bv4Se7+jgpPq1Tkp+H1lslHuRzpjND5ubemT6nf1dDp9suXb7ZUjMA/ulAQMsbPLsb4jH3
jGP8EfZgoBschHnfzH7SoTMm2pcD6m4NuGjNDmaTJAHAmpZkLS6TOGetp96QfURIAGIepP3RSRRM
K7Jeeu9puoXdaVZ25WRds7gLfceQta53N6hMwiTFpYMdiC15dMruT30+3ZGCJgQxjMlpD2JXNMqJ
6ESFkZptHOWwB5AMcax6Ihmi1lkG07nfDP4QDdkBrpRW/jlI7YGQDlzv8JP+/P+E7tyVkr05wbnW
jMAvJcSGEp37JyZp/nJl06PSzYW0PXHr4+7i0pDO7qhU5oEJ87FE29XvQUULgKYBnBRQ/qciNyBO
DWe48Yof154QfW/vLUfZrmYfKmXrNO06qvR18NSZD7BYWOD+uGs5n+EI1s04ExdWjccJEqtRUTJC
nLsAw/hf5/oBEk1JoM5gFsAHbIpSLcPL/pejUVlI38gc3MGFzZhUk9yPepZjdfGPF7iKb81UJLVv
mWpt0qCxEQ9dbxARtinbUBQjPAoBDH9hQNib+iNRKKy7t1xxrSN5PD2WkabjSaCMo840bh0gB/o4
zr5QD8vnnIj6uTqECQcXlZt7SdAPiQKuUDllOEe/fImSdyCETQoziQcwsQ1DH4F7H/lCpO22Gbpb
Sm/X/Dm5JXyOx9W/Qn8z7G3jjs/3i/BvpjeVP00m4WFbfFosLIbaTJdyVH+pIhkdqFjRcNkdVlnZ
HHZdBJJgt4ZF2CV5tuErb31f+vYglp9WJU8WVgqimbmprn/KhAY04At/EK+tlPVsgdEl9uttjxCg
iEeyYGsfU2nz3NSNwJrQKaVEYXk7HozsK+tNSfWPjBh0KGt42o5UyGPf2cVTz73ZbEWZ2HDqwBBg
TC2e2isQcRtlT90X1FPGDCkkOrSTxv0rph9tvMHDplA6dZHxz+VG18GnpP7skZCwop3LZPCJOLbt
ge5/i/5vCqvdROQfL2KNNdr0pxV4luM4xgj0V6ZJsU55B1+bn1yQsRKCePWBFvzm1hG6CNLs28/3
XpmRU9LdHuRKnOavrU0gY7Q4cY7MDK42RFIuWX/wABDCWo1MHA+FJncxc2qGF3stX5kLm4dBzZJ7
FqOqbe4M+FNmzB2U1G1fcU4m2Nh9y4QNxGbSAtMPQGiddF1YXFOwaW1BxwWAt25DoDbHgfFC16g3
sL/h8kZOlXvO8Lyz3F4ykD48uM8nxJDNcgG6Sh27EsbCKUbQQKYbF+P2WPwtE779A/gqD6FMxIzj
nrA/kPA2Zo7kNlEy0305XXz/9M//fPtdIKhGDBGQglZH9FETed2xRAEbrkSDAHTj+JhLC7ggkbf2
Dh3MMnUv+pmf4YDLBK2euaVsuP/gVD0i4mW/AA/NCoPARx5M/sGm7KwXxetAYRm6HEHrqWBTDOd9
qhplrhsFJzthiPnbUpDtgu05IdLQV68MjIF/WSvKBmOFK4ZEP8iHuxuXC89Rg6Jpb596bUKBSxsG
yvG7CwF0J2uHK/UPMLWR8I7r1BwQXu1ntbtpSQyOc1O9qPd8t98xgZc7dBz8j9tesDFts4hNVcwr
2KS06vaHprDmWjqm1rQRrvG21YF0khZZ9TuAGih+mMpjk7c5AStojpo42h+/HIKnA9g28RjeJXx5
sCqugJm41GxKnYgUv/nHNkAfBY65PqlesZvx1RdDvF5/q3BZdsep5q3WaDyXg4ET5Tfkr8blHMqg
7Bfh2q94T+9/czFPQeaTsBITrU9GqWw1zSgttkaTKYSJXauj8QM8DviqAic0Uyt189vgcMcsqwgH
6/V/bUjsegOGzGIk1S92uPSd3Vj4bntETurz5Ez2jBIrO20Dj0ejuxSNIus+1A/vzEzWEonzokag
wG63HwVuhIVdmpajSkdEJKQPwLQ2bVQVzpOs0vkkTfQRq+JX43Fgwajmzkhgng2YjHrJA/UZfWKm
HrcpIDndEYb/7zNtzG7xsOx0nyxz91H5G/zB7eDwl+PE9S8yCpA0dXoZ39wck1DKmfTzrVUB23CC
yQqiokYCIiCGAP9vYP7EVYUF7OKkHRlfQf1B+tW9PowmNGioGqMsHbcSRdE0zELKNx4FXrde4/ic
N7JUxrDZZ0bQTazAWIY/UyCM6AqyInT/Fv175gqvwyk/7UAHaPbqt627BwbHqGhbktwL6lyemSa7
omIk/SsqDaain08WmDEK7Wve6tjKlSjMepdufK9toS7ghzA9PjuxipyQqbXfxakPjAHnKVYzUvPT
7JG81FTavDwmJ97OwWkT1nfaVLHhwsjzVkjMA58raMM0I1NrKxxBjRjR86qxgvHT1SKXbu+Q/ZTi
w22FUxD7n6NyAQJr1kjVJKDKEkj0Ig1ZEbhPSBraRedt6C8IczlBX/6kREHtbhDys1DJtjGO2orW
0fNeZceh6OQGIc4raRVjhAM3q5WlMViylc20K0PeSqKDhOt0LByNbp5AthIr/roNC+a8kPfmRHI5
5aZ3ycxhdZANatB3oTfB1keaSP838UxnAeK4AjGnEA7i1g1HQK8VDH8WP90uRtBzcjpfLZUQSFIV
opwSsfh/sgardNOn5ZgEPnHxEqsmZRGRJseQorC+lGWetjN1GKzxrLmtgCElWWsUwMeNfulnut6K
41burhdhKpA3bSr5DN4KBdkq/OFgzbsdJR5V3UmYUhu8cTWv4h6q4Ha0xE1sSGQN9TXTY8mIcY8L
wHQXTMiAw98UWCN+7fsoYjX4BBnL1AEtReCd1OrJ5ZGH8sbikR+98MOi+BuWT45cqBovx+2rzoJb
n6QTPmAYH686afOXv4KnigPFQ1IhXSk7JKpga4T/ZbQvyqipbUWLfy3VlU7x9+8T1/JLVhtruoVD
mA0EbcvTXZMcdE7xFWk/6k8WiB/aK+UaMiJwDcuS/9Klqj5kpFPuJv+YyOihGv0fYGx0Ki3Xm+AA
3AV/aOFwSce6g68QsmdYVIX6tDmdQtnmeKB+vE8ymTJ1Y5N8dIWgGeSk+C1nNwqXPfYtIJloFfYP
/6HT16egSc42RSpaJdSlf+CuvDcfXSNEo5QboeJnbOJbwjNXNrAG44BncGORCKwpYdHx5g3FEocO
+vA+UCnWuMqkfA4N9iMOb1WGFazDv9TAOkqsIGMsXjM61dCq8+ic2R2g6u9u5k5JztYWHu7OW5ri
EZkdycK+Kr2bMxjhbfBAqIGDXp26W8cLV1XRfz1xXIywiEnHHt2mokhjTDrFIfXm8gSgAwuwBBQf
DTzAgYrQwMCC/d3YE4C1scEArKBSfDg5nRGcPf533HEIqJ97B6VAQIL9v+tF6MnNDpGYVdHigJIH
K4vzK2FqePelX3dAOYBqKusmFnT2VzacCx6hZQXGVfojyQIzriMpn1jaZuN7r1FWOttaIOp8mCUl
kadj7ShOIQKn3La1coeD0I/ts9Y7BMkcV4yhvmhIa0MeshCGFli15Iy0WzihcdlGAqIz79pI5PiK
1rym/pUQMhexObxUBeWG5T8g1f8IW7Wl0raro9bukfjhs3j1hRgPMlCh7MhE5q0koGjPofYjLmbT
6iU8KPsF9VSCJ17jtmmJenDkDuL4UbHpwxoGr7Qh0+0e/flqtOhEBc/bsVRapLgISNoI27vkfVB/
/e7D4/7M+fNDPwKm6cMMisN/xg9IXFe1jn0BjrmTHsYR4uqk3pWjmQE7OgVnaSVVvrfZX84cbHpw
gLzNWcqkfQVJR2o0bspCGCnnNp9wKKVy0Wt63ic32zi1kzoSHhDufbG8/iQjE1M8CkXxPwV+T8oG
gOUUR/3ynkt128GJI2HDkaW3HdeoL0oLHb81qlsOQNyJFv1PckohjqePFMqJNMuHfzMgjcoXPxCO
rSXpNAbdnkeOZ/CWGO1ObLAoGzhB4xL0D4+vAo6aXsjIRVLOAyO5bUo2jg3AdXK7Mysov84VteuY
pa613Dl6PY8+knPutfYCbkXqmYcBq6NSt3saBfg6hxXxQYif8gN/tHQ/roNDdMTSeEcksPHyCvyt
0trPSo1VNoqxdeGAzJAmsz+zOHxlF9wUDqXYxoYRkoEAqpJMsRyuoj8m6PYoeC2X1dRiVPeuMVzX
9yXvIloRI0xQO6fzTbN1owtq6icnu8FlrD5LN2woeBKHM5m1QA+uah6aJp19Nv98hEMEuBylheqr
aK4G4ScLVJrTNrZSNHnPBOHs/0UNzVdTeBBq0EGFJhRThnbb7UVrsS1GtACuQbv22qcAEKwiLycz
U7hkVqhXE2Q3hjoJoM97vYd6s4OsnM1iIh3PjYsrs3raOlbnxFrCmgMJfTm6T66XWESBsvn556VX
soECc6ZpQL4Ghmsm0VFiGC8+Wt88mN8oIgotPZ34+hjHOXav22hrdMrrwScM625RQOGTSEQB+Faw
znbWafGVoRV4f8RQQfql7x+VW24q3ac6t872e475iLk6HCpnegLjzjvgPp4ReiROo9jLO6GDV9U6
Ez3E9XASilVs3PWDFb8swZMd1CGeHKGFKgn+ARzxnQnSNWhv7uX/2XnSHWJ+kWr4CD2d0+Lhvibk
MKGBNqYJIewaSAkgqA0AlcRiTvK7FYLB6Di8dY7794E5cNcEtiOwdr2TTHyDEim1wiQWZC9zPcCO
e0TcLmXA7NPZMVy16nVNqvU9KCmWbmJQRmLaGyZDiQLdahRBa2VjgnkA/oGJRtDQbKDA3D+ahvHE
8OaRWP3qEfzfGbN1wE+8TW2QV4mszBM4a6dv6Nu/GHCXBuH1J2EE/W/DfyMTu6nrKHUglVFq9lSz
Uxv77msjlukYZ7VzCqIQVuabUpFswDT1/Y3thYmRls1xP2HbVQqenaEw01yLZ+dN2MHnF0bV4MFf
qW3a/U5hLHiEvpe6ntr0iBXMEdkl7D7TOzHnK1WiqjrLwv2Gpo0MkqbO8Ae7qRlTg5SdEsQ1SOWw
jtodJVqtb456zGED+5uY+yZKGIoa9qLAYfxA+xdJySm5puzTCrJr9kQaJZBcTSdHLwo6/S/1I5NT
q21lJSqc+C51fbI2AGGxnYyAZdPdDWNL8xLN9V0TcQkorOQLZdyUES871mizNaWIT8J8KEtXKkzb
XhpgLKwZzoSSkHwOQXkjBg0o8UCjbS65iYhdBaOOjoVve0aH38R3BHCu4kxT8T59ZIwIcof5bkTy
v1JuM6kW2QVaTDeOmOzOWdAcIksSrYsTpYta3LMQ/C4Fkgq5cbP0ftkG7IN5s5rJJHsDoDfrUdkb
GF8H5+TX6exkJd2a9DXAdGvkyRlwskvsvGZE8G8XBOA86CsGjGA/NkV5sRERXDAp2qLyzmodfU/Y
gUDlWwre1dXeI0/3q2qK4nguO31l9HcBfS/dmlE6Mj5tr3qYhbx23EdFTT0y3QZZGCZaIG6wuFIS
90YGxI8etsDO6wO61Xdm/uO8devc5cEq8YDV9GMut+Ry1SadBHOci+CMPqXyhJxoBTdDys+5iAFV
BWba6QiW1Whp7KOUAmFAE1ntShPUjkr9e0ppyJgpm62toXYtDSvD2dDg+IED98t0qClEF092/bhW
KuP61e/8grH2260FgFPePk60OR/AodHt1eVvSt5kchQHJmHg3a5vBgYRJQPbO9phojNNhV9MQNIr
u9+Jsf/S9gplBdOJemJY1YQdR5wBYuyD1qTDiUkBzYLmJFT7Bsye9O+d/GpO3y1o6kXktK379eep
yHB7usfiS9UeGMcSi/jf8hP24tkvAYesgFH0ibwJy6tonoPrY0gBZxHZyaXhXlSX4t7LVW9nWjSV
VB/EpmDkTfmWvW3BEsjZdw8ZBwunlTEOM06RVCoU/0BuTP7VZwdAqgodl4cdPLGOtAHZxzZFsomn
Cz+lsQB0EeSf22AQTITO3qtaTnFP7k9B18TWolch/YkGMzDYRvpVBFPMK4NZPYmdTIy5MEzMjHut
PaEBWvmro2EEcQDNCXIxuUSEYcbbN9WbhRgHKC1/9X3NwVNoWnwBr2sQm9OafGpP1ZNY9SeHurgU
6SPDV+PbernEdeACZ+X0r6yr9jfDw7gNJUVIkpmOgIS8F/FSX418ACabil2oZv9m5BIr2WCR+5zn
k0iAWzvlJLd6ChjxoMJJLhAsoIKaTOTbsd6w6EtYwiXxDGYTpoCe/zuPY8VmAElHODFyeu6KB7aZ
9LOhMMtOZaWITUQDjnpqBJALpH1nRL8XaVFKw3cWP9EWgNDKZxjL4E98pVr4C8l266HuC+dfNvTd
PI6m6B9UOLsWXhrVQEMdGD5D9yUmmntUmoCT8UtfD78WF9BcZvMo2MyzFQCOsbyEqY5CHcimEDyh
ofaKwMPSlmtuoBhsHrcRlJQliukLK//S95sAirvHCUbE/oDk7UHwUUUKVhGYJbfQAWvSNPF/fuJZ
vMaH1L9Dyw+d9FLD0rcFP1riyvHv+Qu6UKR4qGYSNK28UcXJG5PpL+vZjm/kCNto4u/xwnDPIm7Q
F+OaSKOaXIGvnpYZBeM2EtJ+FJQyIsq7KCE3GJYOofok4haPcjnvu8Kcteu/dOx1TG/toKM31TKp
vCoqDZ2hm0BBP4cXehSmfPeYL0SXVTuh8aGEzzLvZoPVluaA8K+DEmAcFc5akMezXtMPqS2uR0bD
lh7m6Y/lfg7TPFFuhhD4H/kyGyKIE2l9+dymv39K9HIgI3WM4dZC6j9uF1ISQmEUipAxMfCkYu30
uvcqHdpSvw6SyJwZYFjJHlCaSaIKNBfjqdQ0+nc6KOnNBWYCqKnCQufkEGW3WO8ZEeq0TL2Qryh0
UJ70jWughe9AYhCcFuqKisWJI4jdJolsXAj7+d3LF6oOIocfyjfyG+Cu+b/7+KZR04WFAB5gf5Uz
MOlyiaj8q7bkOcbSr7nfmTytBWHWChftB0JnLKhkoVnUdi1AJreMoKoZ5T659zPTJRoVi7Vy21EL
683G1zpdX+yb36CfNF6lYn0FD/hiBuLrWImclumyO6yxAFPu+zdXR1l5NR0LJbovF63c02XGOGff
ICykaCEYQTSMU1NoTXNJQoDppkMfEj82A/IJqNUXcb535EIZqCMmRuuX4A7OMkFYipL1lVyw9ojW
r5a14iDB64zhIaFkXg6uQ8+XiNXgAuy0NMEMrb/CJY37pWeF7tJiVNKUmgsPP3t0PsLLA2DxyVbi
rOdjDvsMNf25QF1exUMz9+QaSbrE51T/Q0hTz0BA2+c7nAmffwPoYQrwUG6iaJsgVsuto8UAUA5B
GMkEef8yqWMdd59k9GB6cfhra21UosS5PwQnfFWtwrv+PpGnilQjgWsRCoLjUTRI/JjBQ8KNytFY
3ou4O169cFWDpB4fGCoWDQzhdW11VifneDcVdnj2U180hfj/DXyKGEr0eHZDfcYmn9WDpk+307UN
JR2uPjlHtDJLxjzqra4fK2xlDzVeK/a7YUIVt6pz/0nLA34t8IZpnGT4AxRco55SqiIAsvnx34YM
QpxI7FbP4MqPHLfGgsy5fYZIBIVOJj6X8ukNFrdY+LLbploZUMDcJDNlywe402YmkmYdJakyb8Xt
Sdt7zOL+JUDvhzvKbv7AN/u8GJoAIrKrcpNYkUzpMKXqh2V7OI70T+1TXlOG00A2JJWdZOaCwxOX
Yt1OgYlVTt2LJPLtS9LqdfYPP9M51jGu3WDhZhHPbucrbykEPhQhKmla/aVmfU7TV2arRPNM9lmm
bSg0LGUfWra5tx4lJoZst8zBpMELbg5fwBYURuDklkBKekLbe5t+H5oEYEuVrElhuALFfOT04OCr
S7dLoJZaM/kk66emRLJHDNsIw1sR8xiYWESXLxaSNuZSe2D7FqKNfi3jXlS30jeuK7zd6X5h6k9c
dwMfPu7u7LolagcxAT0WgbdWfRM1RU77G8EkI3NgNfZYUPTCklVoZQFWuVO+NT/uj1Dgt78CHU9L
AgZqpIDwuHOGlxvstvdkOTWnu4eAiWTvcCBjz6OAKHTon5Iqoq9sNUfZ2TeZax91/lAVevqyFtKV
Os4cXbELa84jBeZjTb8oodC1QKMG8EmiejzYZXmzzvsfjJwlIEX1buyPxoxTbR0UKVY3PHcO+MQ+
QnYpmcU06iejCvam4FFDz/w4+hJo6AvAwFVn99qomncrsmvRK96QIZwVIaS5sGUsMGfomhuFJ0EX
e4TCxXSLjPBR/n4vaxxLHeWqICQQYVssLElQ742xOaX5Jornj8sQ6Uu6ScRNvMfi8+8lREYorLLe
CDrO9BhdYT8zPXggSQofSkdM5sC6vWxKb4qs6tEOHh8EVpGanVOdbKYOUsJBKZJv04E1X828l2iZ
1wPmoWbvSUx8qE5TztbL8diOBc1ReaNlQoVYMEgN0mxpfyl8smH7xrcK98LcI17lMnxmnpUmOBiA
NcJgx/sIpQ/whSvx2kKXFYfcey+vNQLTLM8pfiqSYtDTxeZv94mKru2W3qguZ5p12iU+z9Kx177u
6ln70GB+EiZ8W+DVZyQJQssl4o8POrMrPhwE/LPhnTT3LMyLuhVuLPbFNmUO9eDq143tVxFhI2/+
Gwl2a6zwHKg0lmHOBt5XdpqKNww64p1fTDgDGsVg8dj07zo2dDFJa1ArPLJa6A8FcrqO6ao2A7rS
DASPgRtzyzx9laU+dsTt6O24Ox9+4MJ83DSiGUZtFy1v3DAik3mz70oMdSuyY4U58EmI7yskh5Y8
A+A2Bn+Zk6zA03Sn70dqtoCpCcJHZmzEiBCy9p2xikkUCQFekYrLZHor+UQ/WsdlCniroM0Yf4on
GwdJkETAW9gjs5BwHi/dUabxGhROzfxHMXP7zED+BrJePjlEDU8vTT4wipvEwhbPuvJx3N4AkEGm
I6ArQeTI1xmR+a5y5Q+eQy2ZCsGhFvUM4RroKWv+DZkNm5UaueHmNm5HntbimJOnASt8ymH1+3Td
OJoI1elanKCtXGipX0G09sIPbT3YSXgtuzvUmP1XJCawYJZbEkd6ResTM7JqhtnEOY0+Pj04kNPN
NYbcxhVTF/mVGajoGRddXmtD7dvwohJGHkZoE1XDugFjyZWesPaE0697KbN/Sk7RA9sxDfH8d0qy
OskFUomnG/rKZ5AYlSxdDjlGsE6DB6LktNJrLhR8SuqJgmY1HamTnW+ubZboLiPLkwIaKmcLAxun
Uho9IDsNBUdIx77XsvNKJ+wNqRNI3BIh+xga4tDt7O+TIVLEHl5maSkvWE0fbrMEjTaYjgBZs1L6
xpHUR3TyIjq8Uws5TJzxEXKOW7A61ulRtjZHEYj86hhXrCvL7lECF3iRkX8HjLMB8toFG7Mh0ykR
y/qgtC0r8ibaJwnPgi/EE+YPbdCXHYsALdJ+BANg0vJlQu6E0YuPJosdOCzExD02GXuHjW0pfcM5
LRWY1dcH7THexaLsTiShe3Qn2wqBDJsYRwk82cZ6bF8BGqxm2KdQiWYVs1Z4rxvHEErCEb+H15rQ
dtczspwjbFzawehhnRdS9qhPU6jDVnIxP3FwZkPM0YjgbC+jzQ0P0OTleInDSr8Lz8wpXjhFqs4r
wdfqsHfOUuvm3u0m/aBYibreFTprEwEpdxv7eaXQFd4TODwpBtUjw5pAaovCl8+dobRyV1zTCNbH
P1+3YOzXDOqMpua8HUrCeb/v/MTJA27xNMINlVNzk/achIDV277UjO7yshbQoZNTgFwemNM7/hqw
jIjqSyGIxEcRopsVC2esTSOPFj8+vLrnKYYhPGHqpdWEt4doOs/NdUIuxHfoFoRYgaZPpiiH0/gO
iLD5RthdywlMLzw9x2DkZjMgomhS+VJw8LbXKHOlmjOlVWy3Cgbmndj3vhuypIENeH0pE6fd4bHt
HEtA+8D7/+EAhXQxFTOBQJ0EVRv+0TLqgqwVFX5fy9vKYTZZN+a3i5i99r8/HTmJiBDT2xYQqc/A
a/VpcHiaO3vLoUYK2oACtcGfK+ICBgkvt/FG6JqztH/jqeIYnTgbYRiRzbi4EiKtPltK7vG4nhqA
u1KEE9ZAGk0RmPtKAq2l5dnbzlDATx6Zrd5+bDgtH1M/jRDg9QmFQ4cTzl5NreQ8YwQMNklSJ7+5
/bIxu2rXToqa9m7MOMgiPa4WJfXvCZO0pv3aCeFnXhX3h4uB6myEO95vXkxIcvus5Vtlvh0d9oF6
EjD3h1jiKu4DRkHWtKFWf2kUkAqDWAW7PmNytJT2qtRvEIC2WHWwqN0+BR3OhZgIajptYPlh/o/E
3Qtd9CdOCPloHBpydghpIQ3XubFRplqXbT+FK5duNZj20m2YBFsxKD+ZRYYQaDtwuRkq5hMFz/Tp
PzLI1Ce0fC3CXnT3WlQ+KL57e4OW86BVEMwEwjyaYTk/nfwPK9FRk5cztUdJ4RTeMRHWnE/95wuu
K54MVEIexRnljp+yvnpZzWLL6ggI+yj4NMuMiYShmRkFudN3tEimAjGqjQWY0RBrbMDTsBe3slZ+
sLhwIRX15CLWdh0MK7///vX2sJ+33cmbD40WB96FQUP8Q1H9+xfM3Kx0O3sQTLduq4hP4x6+/9en
F43MKbr0HTO22TVAUH/SeLe7Me4EXOUX7+XUV28Oci0v5Lbz4+q5COrG8LIQ5DSJhVFpSCGOkLQI
UWqWUYjp2MXUziAVdvpeL+CvRgul/V8QrPkA8AgkFMTtMaukH2d/hO1mqhWuLJ1bts7ScDkaQ3Ao
88Ddf0nL0o+FGFgkGibas3Xa6RZxxtD2PlIUbt6ty67Ko1LCTbgj0n0FisJGkvQ17mmc5rs77ENd
U7V5H+W4aWWRgEsXawFjl0L2l9cVvdGGQD4bg5DmKYinelE/1S6kTdKPeQlvmktuG3FCZ0TddrOw
z7Gq7kmgc3oywjHPJVAsYbhXa0ElME933GGWmSDgFojKcNC8KTksOl1pKXMJa5s+KMk2IRXFkLNM
Kecc8OFfhblmFHHaRhJGjmcZplnNyinVOYAgqrhDiWZm8/cSeKVVJr8PXKtbe7D43XpZmPgenPvM
WGb6gzmHiRaQk014LHi9WeZOeqqkDgKCedeXpFdEWMA0aD5FYIP0Sc5ccUTP+5RY5yixydmj+TMo
yLvCRubncpowMhSxwHc8P/RIvuMQO10dNmEiliPQOkpbWfhWSLvqN5BFBgQh+5rfnH2zzzl1z/U8
1Qq1P4VWwm8NL8gkhVujZaxvl4YZ0zhpUQFUZIw+1VKDwclZGev+kJXFchVPr4t/9DTfXDEyKv82
Y8/IbwFDVkruGtHVUYuZQTaK6yHwZa49z3v3wlJUi/AE5ABEj7SPHttekZl7W9PboLHfiIObBIL4
hrw7Klo58yW453FOFInGA9rDmDdH1SHVfxlRLFNz6rpB60Fe+qYnIacy2heKuGHXbDLeBscOZlli
dT//ELPx5mjedtFCNF1E2ABR1XuphB4vmtRbmR/Md9N2lZrZJqQGmm2eyDLST/Zcak3Fw/oDX+MI
qcO7hiC9nYNhVJ4tPk9f5QSlRwpLb1Kdffhb7wxZVErWylhRyLkXn/2wVWwBEGUa5ZFMlHuWMBNT
ZpEO141qL40wGwvDA11EXZ3ezQ+yPVOTT1WqsfBFzDkLTHNd2fM5W0Ti6WSMyaEOtlM84zNJXcjo
B4fl2/LF4LloVklVERO/z1iiDZQiMpz5lFUZ3qH+tGFde6cgzdhnUUAO6/LanJSuQgQUo3OAkBEg
evbERbdzmk23wnaDaSj1XgV4f5khrhLxkjdLMeToRjnXgZ0DuvXWXnK8oJxAZ5Wrxh/6fGy8vj9v
4ygb68+EXn4sYQlXS56NCoF9/7DqHAlWhT360Lky2c4n/6waowQmPdbMXux4/MxdTspnq8UjRs9v
w0ci1jqKraLs1sbioWXgyunR6Zs7KcXAfl4KafRjEt/u5l3+PueghvN03oWJHcxYN2hkWb7tNB6j
+DDJtsT+IhWCjC09iN9TWBp31jMoJHfKE8qHqQyf+BqG2/Sz5Ur+xtKEVK1hEe08wAeYt7yE+Fp9
SQd25jf/0sbWfN67bCJxRMwnHA7Li96qnIsrpZYA7YYj0+A7Mepabsj4RkaiRqgcVTruuqNF2qzO
5r4nT7BSUXLmd+tSYAN8kUfWe+LBOf+hKp1xkJjeIt1lfyKx7HRXnOcVnG2XJqdVMaVkOXWAdc1k
hOTwwfR18iegtV85QPzK239er7BoJFc733+PzvIVU/tESVMisdoVw6qSqUxPsFoxSY/XhBjI+ZCN
FYw8smE9NdZG7Xd2F8bVN2PgpQ8syGOTfpwDlykmmr3UT2mr376c2IQClDarTb6axOban+qmF3ew
pSXtwGCF+vOaaEnrdJRB7atTlH7utmPvrC5G/Qxk+/XwrULN08lZsLBcXKYJoicCUNwFOsKd1dGX
iBtxZvtYzKcKZuPj0wzEzOPMyD0q0jGYrLc/0JjOks5sxlcTlyulT9Koqh0esuW7hibQ/XzwfrR5
xoct9H2xLoa7ayjWfDOjNflDXn0py0OAnN4KlPlROfEBLoLs6x+1e5HsbJ2Gigko7vke78cokRnY
21oKbJ4S+opf75JTVIep/G+uAcDxwzxlQu7zi2tPPGpWAMSR1TgZc4oAjJrjCjRQsSfI/SZjAQsQ
JRQ8b3Ay0Ot2vUFmh14FSiqAm9/L0eWZgVzoMhjqzjcluuczUbx32aOEy4SM/ZRZPvTVMU+uqZ6B
loLXS8TpSEEdvmUXf6Dhfe+0tvZqVX/VhSPQVchPPYDP8sC2ARrZXPC7JuIbZA1aI9luRyZGB1+o
yINI32q407eC/P1lumB8Qw6UDx4UQTdWJiKzGnz8O1Ed6418zVEXfQYEwx5mhtmwaPuydJZETVPY
Ruj+Jq1LYTNGewW5803GpehkiTZKUcB072DW1MjXm3AvycOrbHa22aYk5nhV9DrT0nq4GVojivDM
w4tW0kWcBB2n9z7Ww5NpgKOgJFPqe/6Wk4wIt2gu6oZiroynUBUKT+r572W7+VtZ4Sl5XXROwP5i
yTkJSrYVsASS8mHIhbPdthIkDjVkXC6H07b44cVbIimhyqxqgFyuqZqu2L1aHfrmi4M/aAp7zZRc
u5xIXx40h7d301mGcawk0CkU6Vak85IvvYpypQYc+L3TP6/YNgvONMEf8vLjabxOvVIHLhRYtzkz
vpjplyvvirUZXFd5D7lxI8IfW0wnuRRe86Bs/m+9wrbvICkB8C1XuPz9Fz0ExiHBZ1HoqVZ9F+1e
DQyR5holCBOA7fHwTZ4UbzWqYuGof0ILD+rf8E52LUwutpnLhXrNXDJVFyPWhhNZxkQXGPpFTWRI
YAGbzLUr3oe+RHmQ+yOTGv3S18onIU11bkZNlTwkp2ir7btpHM8R/HZzIGzWg/9J7Q+gZ+W+VN3g
DIk7YxDoqsbO5SLKvVH/BjJ9vfO6saaoSiTEbVC6yIYNKg2LlPMDwvHgkIgPRZfP/nQD2y5wbEZQ
g/VMJrCnjW8ZiZs7AagfsROCIDeLwCcmKvEfv2f+qaZrQOcEGs9PVx/uqsYBdaS/fNfUdberT5jc
l07OQOMjsUL/8VS80eI8Lb216sqkxkjqq5sUTqdinv33XQgg5/PZQX6/wcflfMvdsMWzpQgPW+Ys
fgKYvJhDU4u7tAVolq8o3uXQZ+pC7Bq0fmQBfooSPkgA3AN9Uai5VUl21lRtBsnwLEtMOKQVEi2Y
PMcX5ndVUDNHcqUBGxv99jHnT9BW1st3rdXafvq3WXaRLlnvSFivjteCDxLrjTcRtlVKtZ+Mfz0l
6dae4niYBV5AiOzVBw9rd4Nyg2yMLEU61eYmRXgh3jJZYsEkV3LzE+S7ty0+GxKpgK+7QqG5DAV0
CNJcNU28kbr+URwho3FKkCiF4V8bq0vm/Hwe0lCMxAZinTWST+IVEfoAoDHvYeg4Ow3eXkSlFwkf
nn0+uVU4KCOYHWY8iyG/xL6OJWRqzdEOOdALZ+OCCXFvz6nmtB3ipTyD4jnuJ1hdz6H3uy2xHW92
BMea9fotxuoSoRZAvnnR6hmbiyWI4UKurcIQ63BrhjICXWfDk2RgCp64Bpaov4KX+K1UECU1yFwr
F5x46W5irpocm8x+5/WBcdSNZNPOOZDwDjoylTTiiXjEsI99782idpu17BzhVxWo8tYfF/FF9vEd
7BrEIMx/JBZOBKvi/OVeA/z7hb5BZVyd+iu1ZxAFPGFcaXCnMnVIWifqnhXm1+S+FUkmz3lzR2Hd
YkFRac0usruH4s/W3WiuZGutj81yfdZz/wr5dVybl7G+/j5u6ChQOACXvM6pgZTLS9CGwjOYtSBC
3j/sO/LjtZcMIMhiTTWg9antVGRsc18wZBqyVkd6tfPsL03UQqjzkwAYcs7l8HrGz9YuBQpGhOP/
+MQkNDcHYWNhh+BfLMUfSTdnrjDx8Cs2qaGOEuzB1vtUDiMa2TKkWbc7e2eXnFvc6izIQ93W5K79
4+uFa47v5cfapZbOYuA0PnMBw83vFoX6ATlNtlQUHE9xTtC+T+3E8DmSPvr0zG+5SeU3WsmvQYQ+
4cSPA3NSEPhyi5wx4OmVVnJTIo6mNV0X9maCla5BUYTS5XRha2DTu6AjAM8i95kjV/1dDhbEUFxb
pbd5kpGGQsXf95+L3HE36diApz4CzaONJ58F2yxncShHfpBhibUBHf1yMyzwQA3tltWctaa5vsHl
w/umFinFOcEuxrxg4ulbd9Z9GSwHwc2anFa+KuY0POZzPo8NPgqSzvz7YemyFyAiaA4KJIQWdhZh
Smp1DSnghRwAJ0jMWvHyQ/lpJwFEn7uu77skzAXPby+SQdvHJlbtWSvRyKmTzLEkJ+9lXar+Bc8a
BVl6F6W51ZlW/aWNgcIgsz+NszTX3IniSizeNOa58QS/pE78egg6jGV8ZyKW4N5rB0MWLLPWB+LT
eKbRBLVIrOwhKQO5ylemo94OxIB/GGepSfK5X7lBP+R/b3+ccZLs3ivgqucizX9jr76+VFcOfz3p
HS/DHdTldkshLI2FGV38+M6sM4rafRP7wGZclYNDKB+1GRYsTyNMdn+MIt/LVt1VbJCm08r7/rQV
0K8uxyqcRnxYiF7qeC+x2I3x0TkpZEvpiKw4P0t4SsDcgqX+Fa3yAsusCk2OVrjqEyL73PlHhMEK
olH0OI4yIcV0OdqS0+01dgc1j92Jix9mJ63Z42N2Z9HznvPqO5nvhmuoIBy9uZLW51VVL0rjdX+l
Ul1uYZlpzXYgwvBUO7aiIzzNWn8vqPUEs7Z9tUFUynG+2MbtMlQ8WpJC3TEonkvBF65TCgpCWrs/
JR1D8FMt3j45pcOeltWHDJ34UkoBtNcnBbb8Zp8BJq5FP7mMtmQZncNqzmmVpuH1rqfcfDJh22Xx
EpiH4TCe/9HBsJqrLh/KC2AmzIAX1Kjy+O7mfBRg+NR1EI1NM3Rz3sTyQTbU1q/ua4JX8Gn0bNku
5I9TVqTxuVIt1N1E0yZGqLhdfUZUWiNvnyNHkZ/3BHw49ZJTYqIAHZAQroJLpYGVAjXtRJpJxvZS
sJEDMrr9iBG5NkDM8MaZATMOv+jRuZunjRkeJCL2DGOIPQW4BCtnxygZE0vt8fuFWTvI3NXaYSFA
nJWJs+JmbSJ7cxsdn5x2kGB0v2JBVNS/PSyhFdtbUnX+cyYJ2mdBU/2C+qCeTYvm/YSkgb0JqZSP
pdOaa2gMNO4nRrpolHR6ugde0Aj2pZaxaEWEeqClSb910MCPeR7ApDdgt1yeuR9P/lS/NKp2YVrM
ym37NZv2xzINPV7O+LkFiGAqsmN4jlB45+4c1lLJycw01XukxECRw2Z2AjXknzbaRBuXckOrIhI2
UZiHjRtHA2wH8G4BY7bh0bme5DIrihVmf1PnDU0PSuxyZjkjVqai+nUpSBMtXSHvfYXTQJLzht4y
066F/oGm+3ndVWn9Tdsvv57OVTorKDGvQSre06ndnOa6jRiKPlgnPJDzEdnk/newKgSNt4VGp0tf
TWk+9yQsnTbze9j7Huo9b4zjOwmlA98rP9cL2o4b/w2vQwxCuClRHLVfIQgMjjQQsf4vy4xpCtOy
knNZLAANOm+NAjly8FENDrorLQDYwbUo0lcxB7rb4LXuxrK6p9wFnpZKvhKH4RlJ6wb8BOZNs+UW
FpDFsWPOn6sj5QXv2WfJfY9tYyAX6v45qN2+cnSymijraad/El6B6ssi4Sgzm3vWGOdYyTS4l616
w6HezENSzJl6mRRGvpQcH8OwmjdYS5ee+ETe7MHZXjeJlcRwbCRCsbwtPhhAzutZl+PBjC4QJX1H
ZNvf4xY/VTYNoDMwQMZ5aQH3QqhWTMtE9TdsIZHzju6wQprmFwoCaI21J/CYyM8ry0XFCN8YUl0n
G1XlVdFCme14GZ8Y/N4XtLzSQi4l/fMyVQzPI8KExmBC7WUhqskfSnoMKoS9Qz+6JPxabw1laNZH
bPUn9aEfLBBkpFnmdI/GoCAhiVL5Al/eSXtGrD4e2xmED9VgiPpnS9HyR3iQ8vvS4GXI3iwqt2gr
d5831xG6USeDFfcoTDycu5rXzPFYztbYRzjF7RPJWnxIc5w7A10ad18Uh5efLqqzeFAGV9BuOIuk
tV3T5mLnoT4PPpB4/hbKEKyj8kMxf1XD3En5eZM5j56Pci7ZQdHG+q3cGo3CrW8HbvyOlx/PEkBy
EXL2Obg9oefpZ8cwaMfDkKAjE/HstenYo9bE9i3saB0kgr2oIFv79pkoiY2R4ndldj48IB3hjS8Z
feV/DcSDFJSJpgVfYPNaXcTZ8nPy0HMSepfx0SrZE6sTH7edypN1X1BZk4KWIi2eTWp3W7qSnsfn
pjdCWGnjHhbA674Svyv1hj6DwOPrJ4bthMSecre1O6s7zf1hf1mbh2MJLGAUYiiu0XfPt9v14MFd
tdbA/mspqyPd4t7J9HRhfy57S5Nt19w9nWONgXMFuNtfL4z3/tANCOn5JGdypk0Sb0n3YQecJN9f
L1HeWHua+FV6pzSq0s4InhxSYuYfHLFvJpKZMQyOfiaoKw9s6taOEhwLv1bLm799r//jRpQkBU/r
1JmFR9wE5UyURIEE+in2XPIGNM0rOHv+aTvBv78/LZa0sddWzWeW7vWsdtEhjh7jpXV46/188CsM
IZbGimmoDXKXIYYxxg2zX0I1rkGa6YXkKPHRyJaWinWDmQ7AJ8HJT1BZm55KO1gnsCNBM8Cm3BZG
o9wZ00X3EniKnCLrLJ7utP6kOB06QmwS8jHYgUsH2hnvyJ5dJrAcT3dDkjoHnr22TJ6PPcCc53lw
tKyuHcGHti7F4divsDZ0qkVR8rHFnkUa2+Y35x0t4eK+OMxec1RA9lmPndAI+kr00XsNJZZc2NeX
OlkC87uWFIc86vfV9ch8kLYcC1mu7uS+N2o1wCdf3ABMngZqBvNsCnA+/VXMkl/AsTbROAsvhCrW
pygLOCEt518SXKUlxqJiId2z810P4/2Y0fp6hGHiVXeDvdqXBxM5qKWqXg3opOawZnftTIbFvlC3
6kuXIRVXCHm0CFnEW93uDTZ648FuZYq+NU3j5Q1VJUHIHld2jjbkN2q37jk/7wVc57WnqsCo5Lnw
pBptu/n8+LrJ3N11Tl2RwPwWNAWwQF4Pwtx+Sq4PiO4F0jZBrTTOLP+FdUNPb3CLtXFoqSGuFdtS
ObgTZoGbVIaK9YI+1S+fTKV5oXF18EGp6AdUN7EQMhaI9POoCkY8t+i3evrH9rUJozVCJaAt4dMr
Up2jurlJlAO7jBrm+MQPsW2CIwGoKJDsL4PFS68dxUgV8AYddRKBx3GBx2e+D18UpnSzujqePxfz
R6b7OO+OaQj4hvD0TZSbcM6+qjjjNyF9JfTjGpO0KDzGb2nqQFyb6Jl5cYgHyWBqTaY+XUF8OsKJ
c+DDDBn7PjygXUAC1hiRM1gTBSa8GcLW1InEQI/JUnqKmSrbFko09+BzIpWvfdSoD3jQaXEErMJD
YxlT4ekDcjpYHU5Oi9sIbLusvn91f2yFZcr6a/um0WPy+gcSIyrCsRsvzv79qSSHMHB/hXhg06NO
N0X4bG6J5xaSdlGCGWmJXcqWmoS8+bK4vgil2cUKCHbMPkN3qNjWH+ldULMhJfGy1o6bjV2sf7sC
yPytPXw4ayhExgZ38FtS8LJ7BCdg3qQe4RAiF3a0CHqZR38IU2Q5+ltfvto1WgnDaT5Wl/UDma3g
bVjDw1EEBYSJZ1vmb7lENs2o/YQIOvF/5lVGV+ue06Q8weII5+H/cQRpa2dt4FXTXNBdHv/lSdbx
Sw7C+OJjUiLP6+6gbaHj/onZnzWEGygqvFu4dt27P5nLBwa3eCj6ZTrdWsZ2Do2yxTrSK74r/hOI
Pttfjbg/Q5n/5AmbQ0musTSZwUO1oocNwq1ptkkcWEWnaNXy83t4pfNAtkmgCFzu2aWxlvPvf5kW
J38dVZbsNiaZG72CDJJb6GnBZf7oNE53eJBbeuQdCK0fhlUpxZ0HLdkgB2fsYyONKjkgO6rteE6T
d7Tm+Dtk2db4pfbONCJL2aFh0jwGlSnDgB3prW5MbR9xQPWER+e9mvemcZ+2NbUyoZd7sWq3raRs
ut9xTLcokEeWxZhJlAkSkBclBZnbulIToacaXp9mmI0QOSXyvFaAISWeXBHwI8by4HLZWWcR6iq7
3sdBj82zVMyEgP0V74ZG7E2QUv0ddsEMgaKJ6gJVO4q7APsLInQ2arUlRdQB98WcLUv1+n+Dinsn
5l/Yvet+X966Y2bvBOLTaaA5CnnIGMKjnZtOB8ZiwlMKn5y88e2++YwWVXaO5owBvEroPHMi9QPZ
NshkSlLMl2vwQPQQep/gW0eGNbBfJ74+hvBP2CZQRP2Oa3CXoolt22WWckQ+PjGc2ma4NrpFqc1u
pzvp8HpPvi6752IiRkVSlRu+MHiQ51+pfdQ12ZZU5/u8xTduIgn9pGBHCyC2nyjl6/7Zn4tGUSx7
1iqXnEb3cKFK3jLQkhT3CrSNBb9jwJ3Y1xyPcMqwFxymyRMil0Vx+AJmziJ0o9O/CksKJmbPR4Zl
0kJeVcKsgrtj+j5uFMulx/nI3vfNo3rP+FuzgQMbBdK7nTTMmc9P5TDswU3mBvbwnr+rb9J0o4vx
e4jYNr4vv3DY9JCFbqjnGqTX7TkxETunTVs1HtXrIy6CnDvRGDZFwnYwZ/LL6zMj22ePhll9dRL5
58+CszGQpsYnLJXbqaTwtpwhESIBUSNu6MDBX9KMN5UsTEX2OB3FhzoFQggQts74sEbAZy151UVr
xioXXR09CWvY9RGg2n/dXe/A6uiUTz8Z2hvEwOcUVr8qHFbIDBouM3gm7S4ooq/NKYpcy29L6VY2
cZQBy9MwOUzkSD/UxRW5+TulfwXJydr0TL9pzErXUHtyMU4svkele3RJsda0qjYbozEJiGx01PKy
eVX0zPIf5GeG8wqdgtr5J+LdR+nXh5jRYTFeM3hi+PVxNA3vazRUwjgOmegfNjVTP1mhJ//L7Ed+
1f2WagzhEaaBZTOYk+omCOR9ZKR6QX0A1Ke0IB6QY2xh30rMdAD9b44wzeXJU4YJUJ3ZIboDs0NQ
8gY+LJrRzfqdw8V2YDQblD8ierDL+v7LPu2+fIJeIV864rmAjO7izNio3ipm9VRQuMZHm+zoyFT2
H67e2Ctj3dLF5pQMGOz/lpqtDHp0RAabIQb/o0/ebgOtl7TYk9WxhFg/tZ6OGs7VuvfCp3Sb3Lor
R0uWNPldiRwIureZJTEb0uP3JH03F7jvwkRWNCi4x4yr3r4RfbtN0n+7YSe7bCllb7SaKro+rR22
ueLaOmLgtIqNbNoogRullINeuWvDlXRe6UG2pffSyGtpVTyK8zkEb3Sc7AV750lvd7gZ6y8Cqcf6
v0Cu1hK8viVVkBelhxuI/ZB2cTNhshnLb517dv0r5SGO+EfY4zN9qmwg/h0UsezLTp0lWVRVVdaZ
Cotn1DYhSCbR1FoI1WK32WQjlPRSNseK83+Lup999JlQgS45A55vAjwJmCd2dq6ax7MWAG6vpuou
nD1LYWHEfk36SVSCzx3SdXx0omoh3uq0zciVa3k1j3LOX6mTPzOlRK58bRt29ib+ZcQQ3CQGGHJ2
IhQvD9hZ45LBYt+wnXL2kYbohVe2owpS6aDENGHpN68HB2E3uTEwm9TOma8ywmdfM2sUEKDRpZnM
qiykvEghrfh7PvPLZOvn6w0BXd8Il+iYxMtUUcJB3heGjkrOEbe3+lfElN3bP8qYs4Fq4VIfzbYS
elmJVqYxl9APqZL8qKnRpY63xjhkeXPPzW5tGWhAPQYgJIwQvP/UFo/rAzmfIJyzYA2243OOZ4ty
1FI0zYFIUgAmdDUD1WXbcN6alC4J8NDtKClOXLc6lsNc1/ErTYNeovCslYPvWKrlacvPM3d9nRSY
KtUOrTR3rsi33jmKth4orSP+KkEMTt3UkKjSpQrshd67swHTjea71MNF93g2LnMIUWexfEet8zN6
rCsFOMrUVLS+VVtWfijD3uwyK1XyVfk0pINJ6cX4sZSUOlreELYKTmXfCNMXhdE4RyuFChYQg8T+
3l7+ohb36x4qpDe59f/YNBYQ/C3bSwyZg2Wx3JYFsBKzv/SteKxpbg9BVQBArLzOxFVdsA/gfo8c
YXyn59KFjmZebfZo+Ypeu0WoTw0aw0JwXQZpIB3BVrJ89fdVpN0lbOgiIAZuzf2exq45Db+KD+HM
8lFRzGZffzZHcB5TVqxByzaTl8/fcVWQ1rYBn4xrVYWnZNqgMdAVbT5zPPNLXqjqruSaEzYPUtlB
SIJrFrobm6xsh/gfh3j0SjtZBxihq3kfaBaG2fMwBUTToTcsgMtM4iPoD6YGrRd0LE0khJrEantG
pyD1yAN1XmZRt54HkQE8O0yu/PWW8hxKMZFoTKacIB1D3ylOvRqi4+IHdUkH68a6NGp9LdxIngj+
WxqF/J1I69XKGLbuTmMyI31GJg0krkFY4DDCtIgOXvtTA95O/Dd9Ua+9Z6/yIG+dKMhOnOTx9mL9
DADWKKH9iDzY+sHFCDR14w3AkGUc3DOyolMwLtr4Fgp+atTjSQDmizJpgTuhWfwwyJt37vNYvS8/
kQ8eVLkvcPZOB/XLUUD8rypfkQ/7uNH+jJtDODKmLa5jmBgjmW0cWrtp0+R/fpFbG4JwBC6cRZU8
CE4b+OPkLx+kwPpYCo4ohphdwhdXNavn/aBCX4Gt+iFuZ4MsQMEQTc0cTj7Az9czySEOXmXZihJW
nkHEQbX73nyDPqi6wBqolN7Lx230hJ0d9v/2tMkalXaSHyRYsiVYaZGd7GDTVLaU+EKyT8boPJmp
TNk3VBFfE648Qn3qo3oLQsxJeY17YCHMqOVr/NXQEX4Z+mdwiFmUdD7NV4etTtoVAI7c7DCefrt8
O69nz0Pfu+9ZdlKD11/Abp62JlSYihJ1KbnwBBTSdO1PKTyzgmHz2AoijknVKv8qvLBqfel6J2ig
R7oZYNfseE5O8BF6lgERBBUvDnA7eXF6iUtVCnKSp3xiTOVgZVsn5Io4iOPNk/6ECaEN8JQdworF
DPEZFHl45IJ4AUwIIyg4r5Fzw336mMB/Gv14bdIH0qhdSzdHPGpwYxpHMjkN0LnLLmB1EITF4R7h
FjNaWLxtOBdTzaXLLIN2af9L+ezJVyp3hwoUWErI92foYoG3w4m4avZn9AkJ+Mn3nqJfLnDj3Tk9
f72InKzN0wKg16jitWY845iAbUwo5RKswOWbtxJYlNkMpPsCzcy3jAHQw/mcLdIc/u5DuqlQ93di
7u5B5KCe4AykkQaQJf+g5l0lowJjJVLxRcI3clvJxI9hffDylOsXWRj8CiAV3F0Ri/B+Jne/tFcn
z8NZX5MGQ8ip9nPeTiNNUmiZ1bTk9uSi/cUGHUnzKx0Drk13CKAvwEqGhodHAfZQHakyWEHAPluO
gNZuDn6ernaSlz4npeK3UMKR+Tp/pJ6pfm3jVJPHInlzgm7LK3/1edOSD5hgBhIpCrXXRT6oT7hP
IXUZy3D6GKND5QEKnzU8smjDEKhAeAQZv6t60u9nN2RImlowrqZ2nIRtRm7/WIdvYwNj2mSNWRgX
m0YeDUuHV6OqNb8ArYDB2kyl3RuRrV1NrNRMfvZW/TDo0zxve/5UEcj0SJbs0AQ88ovELm00wHp9
byqK9Z+iRWq7un9qKkRpNPKMNBlCCpUfdOSdQxiw+wT5NysEU0Apx1IOqgFouGCRW/wZlbCtGqd6
wC3rJzfMPxiUqMjLOqLTQyPWapWdJua/SnXLU3T5VJNVH9MZ4OiRMmcDYiY3m1hL13WPVPivdUF3
md+ONhNJjyoZ6qzFhH01hdhRa8w4xyg10PoWSrsmyZnfD6LV+aeRzK9uKB3yWsMghu3zK+ttwODT
w4w7SbYwiwhU52fvtKKXKDTrfjn3za4tLF3woEJewB3lI+uc0GNzANqjLoOeGVhS3gt5/GwnX8jP
atPcrmAHQjyX/iqorNk7183mmA7eoYA36SznVSrQ0fXIfoPkhfHZRkw8GhTvI2aQCL+HwuomrC2o
X3L8x9/sNqBJvK1zuy/wZBb3wW/gLT8/6ioeWpiRu+tSfCK+Kb8XQoAOs+twZ+ca7wrDLtfv0Fhw
+JAFT0i7ZxBpGwtyu3AmKfau7YSvOo3nj1R8XRyryMB/aluNORAri+bIwTnacnjU8kiV6hDvxARK
VGcNtxNnbB9FoXoyDKZ963qRtZuA/RKCBfSzg7mZqKxD2eDHOLxlO41DpHSaEjnHWZPIsDw9eMAa
To50S+Skp2XYQz6UMOCexCB/MLx8w/0JgmJLWrHoBQZFV21EBKSdWOlzlheOkwhpv4CDiBP1IGRT
AjkZ9+/X4uJXV+FjuMWxLTEXAmheQ2HfmWsdnj8yVlvo7m+NJYfAEDeMF2DgWgZNEIlvJhKg7Wsu
XMQTdsaXWetjLgnM2vDYAueoPM/vdjZaMkamCe2OUI4uhzRCEiYP9ay3JK4wHFCLAFaD4ceViZ0m
JGbp8DSa+g0GTXvXzy7Y8+1lRbaHfjY7pROpYhoRFluot6UX9fra23y2ulRk6vrUCsc2OYvz1fOW
dc/0boJBn7CVYvpLReASqxe2wdqOTHdL672q998VY0OjgvOOAP7bAXAwwtjQRxvBnZcskUo4dChC
7Buzt9Myr3nFqGk5Me9Txhg6aI2ZJ+3ufB86TJzDT6ARrjFR6K49LK1eJ/+OsDNn7IuprrbPDhtA
okKcb0y7Mevg38Rzurs+lykRB4UaAUoHSjKN76/9ik0gSlnFwu94eiycfPDLf+alkp2HyAuRmLbb
whVfbicRvFFRT7L7Bhw95jy3N0VO4sqszrT1IBYiBnBeKtHIVDT4CGV8CdIDCdWFSd9rV5nvoDu4
yG78iNYnrV2yTUbt0dloq0R86cTDln3pyGjlHQaVe9WdkV9VROU4chzeylvSiINoh+uQpinNUnm/
OQbdcxDMa9L0m6LDaLQ7x27qVSreuFuJpIViSowx/xrvgbXVlClfRysCtwpDA9GE6QC418Um8rQ1
Su7HmGoLJsJ0INlZkvYbJHEBUzlFKqCEz6Dh/n+TjvjAEJKma1IGkvzw2WBNLz1BdogM1XahVaFU
U3Rg/LMuRMKDivEUeIT5TG475pfGS5p6zD0MAueMpqkWYcWDhPV3v8acjnDNbaP2WDSj9yN5qFzc
CmtDi2V1zb0HHcq61IiTA/M08APoTdcZ48REmN68TnH6xV6aRw7cWFOBB4MxlS67Z2+dfCUPwQ5x
P0ZKME5DNbaXDj8T4mEKgYTLH3yMvHtDwVGCnoERkWbG3XwJX2SNysSYmdJjn3AhtBodYQ8zz6r0
kIPsvtLQbzWsgEj3/P058VDixrwKJ4wQZCX+JFpwa5QiWyF0xDwpTSkYfWtIAyakQe2T/UCYOVAB
WbjWpwUMRDPk7S2HTQ/32ES38yj1iWVpx/X3IzqYOsNq+kzeY1iiv97wBq1w6V5kwuIYDF/kwFyR
ePpP63BXBzeSbWKpKUcqsCXwEO83iiJUJYxtShtVuGsw2Yh5DJRNrCh9b4KUCTU2rZApapfSvfWd
hb+QAi+eUS83iTrfdxO5GGSm4CS+p4bPYJsJ2n0ZtpzmLynACxddiWA7SoMXh9ptDDUnbXUVAJ1D
zf4GdL2rOERLjyBqKl3Zz+4GyG/6gRioSMQGir2dB/PWq166CaPuyFZczESIhkgfevEV1lkLf4c8
vQkkSh9m1Tt2haqnkyCcLNJCvMfFs9hf9arlKiXU/I1BiSvGsrOLWHbsYlvhMKIeH4GlkhLdLWqV
5j2c9I+1aDjfCJOVLCEEhn54C6B4GTU8oVstHVrzSMcnx3JzfFGI3At5CUMQu/4f4SPm7CgpYG7E
SXTeGvF659kOl+xo7iyjM45KlVrcLjmVuVlcLHNEnCldnx3m6QIc+wqBMkElp2VpxC/J2XNBq4co
qQE/mzCYWu+hEirtRccj16C4bxBPgB/s81+kt9+hZ0LYm6T0zjlpvzqbNtBQvKBLZX2LJmwm+pEB
hcICN6VqdTfGO8p9+91UyvFqwMP5vidTuHMxYqQSrWKosSGisW8k8uRlxpWEvD90jhkwWqzH2MWN
8tbqk4L4kBWhKBDVZIdvXHg9d6cM2b0D5etn+nsw0izmh+u8YmVsT4CzeiZJED95v4QxhK6YgGsd
7XdJ52yPO0HtmtgBC655ecr1isOksCtElGPtY3fcqaWgvE4RmXWJ3rsGbG/lHglK98fOBl8d49Qw
7Ls9a/f5AI5P82qXZR8DrKKlX/KQMeEIDw3ADeHg4fq2UUCxdRBYoir5QLTTs4smJ+uCdjxR76lb
pKt//c0e+YdB5XSSUFOnM3IqNSOlmK1aSI8LFTupiUiHe6j7g8zr/WaapIzNiQQq3G8/8chueGoZ
QK7ejXfABKVV3UD37rdo0eO5W0KBIg/vT7CN6hX6z+/5wfPB9umjErKS8jhXMTtlheVWZDFsacZD
LyYQ2OEkGwmF9P8tHPpqCsMoDd9M3ENM/H316nD3PgzcFlZ0785a6y0Vrzs/wK/FDdpOLHa4vipv
dp1qDKNEjUy7cExqAGApwUIB8VtSudni0RXZCCg1R3Bnu71Kg5lex/xX3Fc3YlO58fy9W5p+ItzQ
I2+8SMnK1+PFcfZkfXxoXLKsI59VBRh2jzmdJcNKDwsWEGDbxkV5yuvkgfaimQIGO89hzTJJpvwS
kkNvTUzTbTvoMYRHwBefy6H/XcrgwHxyU4aYZMMrOuPbMpnI/FsrGgErcKa7k9LOUKOKuv1/Byvc
zbHLeWUvfSH7/I0oPO1K9Ps9cM1vygNBoXiKqQhzpG1w1DCBloyeUwTxsaNIeIEXlkUv0pjJnbdp
Iw196YIK9YDq5LeyP9bk32uh+bE0p4jmOiGTdbAxTbZZaNd9g7aN23xGJbGWt+294rGW4C5jxCPk
3dM3xP96kKDHb6Q1stw96xN1M9MOFmT5nclFdO22nOug+FaxnVpWQJ4fke2RqACAkiPpx2jvCKII
NQfuIKdlKCrq33ce0dLtwQFqO8aRx04mqzVvLtuGkGvIeU8hAJsLIapsBCxb/gho8Ygod8IYYqNO
yFD9eZOUp20OYnYyPYhzS5HlKr9NlV4cngaTHnGg8AbjmaTqK8jxFTxFzzkY4xJVd8/6pvzHfHWy
SuOAOFPrMF+QqXvlW4tZZmM4Cwh3QnYkbH9ICJMoiPquLgPJyVXz5W8nHqoC74w+GA72DK+4BDtV
cvpMrbKyfZ5E1eggFayWpM4ChvXqWDc8c9Y1SBTA2/NbRA0ADxx+Sx2uAqQ0ngvlDhYVDkhCogRy
aLVvNSx40qEKfNzc/RlwOKn3hlhq5LXmz7ueMAy+d2la4t+57sbCOdOMMlWjmkrtA4mo1wMtDOPE
4wX4IXWgecYPx7x7haTOxhq9ekt/BFeL8w1/NxcQ6/u4okxfQafqG6VA88Irqg/3/sH7YP1yCRGP
NKdfSvbvZCFBb7Azfdw9HOEjTh7D5kfnHGq7zWYiqwRxMI9ldIXJq+HVe51KqFCf7oDqMen2kIjr
YJXfOkvVfPhDL33SBan1wsf4/BmN40i0p63uE29MVigSoStCsCVk5d6LNAcfwNaDMv0tQtOZa6A4
cc6zEWkSxtudoVeqYggKWc2tf7ltyakJ9YIFvJejuPtHP3ruNKahHc9ULMpDB/bBSdXlLYgpQjMI
nljMynJWJbDVpP0uzKGWBd3XRZESvFX0RuaMH8/Vn370hfiux5OIqwipFENv2pbi0PONplu5RmrD
cvxx8gbGPbdjv0WQFGEOfRhH6xOL6BBGbuMa32SCC8UpQuiYSJX1Yi66+Jadwgd8hhP+qYifpBe8
wvUIq65b4ii3JJFZAj5INcA2Ng82tKt/dXSNzIAg6qj5MIyYFylJptmbLKVMZIm2hTJMFJB0vHWX
k1suDdH3lPP5ErvrMKZEMRs8j/mXaAkNcMfUHnMVLKebo+hB/785eNoGdnZoGQnW2xJpluDj3jbH
cz1I6IxbZLrUZS8eTtPP+cms80eLOw5ODm8faafQYPz14mlAxvunig4hSU2u9bDAslls1sGn7/PJ
r0BptntfmZWjOVuMuWknPj0qbWKBPP296MCDtEzG3U29SOv3bLhPpIc9tRV4pA/LzVAf+st1fQBY
9jYzcdCTHng8XZquxPp2etvFY8ajh3uYE0O3PUwIWzYjDRKSSMisE/uP4Ao6s703GKoTvUXc/3ok
sUQn2KP7JCgO5+KfOLVvilxwTJRL7ya6QSxoth+m5KQ2GQNuk309v7uku6ASJjtVfKmIvbSu4sKv
w//idNYytyJ7gS39N/c/vxy2eIgOcqI8fmuElT8u2vFl0tWblzbtCrTzBXDeLoVZuywIJ3RJADUj
TiYwHr1nXqTDTvCoE6e1yi0gBXaHGZCdVgdikWRCxLoGWZqToPGi5C5rbcvIgYksYW8Bwn5BKKiV
e8Zs4EU4hSrB5UAdJSxkdhQYlItRKeXYaWUlcx+FOvfzjjfaJvbtmerNhpRmtsq+TUanNipuWsF0
//KHPKcNOnJ/hZyCoRW7N0kUyfZF3612BcrLCoaL3u+2vb4mKd0SmXHMv20hECiqtktEi9yn1Beg
l6odbtpVWuU1ZtRRoGha6LhRkz+Wp89nSu7D5trR/+MbHoh1gE/ecw056T/gV8efTjtkPUjxpycS
irtcuL5XmELwTdPPqURef7E9cDQMan6E2CYoNmA39fC6Kwua9E3JZJCHBs1wUP7i5q6wfCUjct3e
/H6skzHgN54qEDUx5K2WBLE+A/yeQz737rgdXqjpgGTGidR5iWzqmS6z9HEJUVt5wdBlUMeD4+Zy
l0YC2BkwkKnhGF1MAA8y5nt7wVdgRh/tLJc+fQ5gXR3h0drz83RN0jZuaNK6vzia764gZ7Tb3Neo
+ehu0a8DK+y9341eQgaM9ujSs6RkTdvx05j+VZtjCVIo/IlfiFqXHCqtOcE4StdB7xEjTzXe6BXJ
RFw4XylYG0zE010eSGChIv89lD6ge2Kt+t/xCrnsH09tm8deVmwkNcA3CHyNdBJuv6Uym2gvIkAF
U257iPECtXvQfsJ9LMIFOntPVQKYaQrvMpUJ9+WWIkK1HqJPorLK8R2aAjeiZe1mlBCYmZmh5ttJ
jttDM7VXtTmyC7a0IbpBcdPOvmm0CII5i9E83XaUeWdHEnj6b64rO8cyTMdxWS+9r8/wSL77e4H1
iLjX34vWimSvbYCvdSFVkiOvVoKz0x9yfbwqXEXtEzgzY990gRooi74MQtNIkfZsNEzJv9ddhcwk
CUKzFCY14f2TyhY3nsjelDgSizFMkI658BObEA3JRqFP06WTNNzQC2KcGV9PLey/2euxkYctl/77
X7mhzQ7Go5APgMHHH9EsvdJWi55OyvDTrDm2NDrH5k5NzBvnMXd/mIQ0g0RxNEyuoRLaqFUehBRa
pz6z3mG0yzWHp5nKiN1n6VTAtSzO7HsOdbv3h8RKyGhgUD3QX0YaXVDLZ2Lw4Y/t7rcDcbPpCZRe
SNFcl6aLeavrAg+Ji8Lpgei2vLG5gTLYrQv5HEteRhMkPScdRlt2E1rEJ9OVWrJyHzE4R6s1zyXF
G72aA3Fq9z1UHUsO7Mm9jUDoQBkULs/p7zWpwsFxkfCiwM/8jcqphqtG+GItAAdRyzh30Cg1QbXI
JWL8xrqI+UDcEC/pvb7ZQzpadTxXxOkVPrtqjWRy/f1CsW1dcROj2dbdgFBZcuBKcE/lRSx3KQJB
S9RSWX9nm0g4ctPZyOpT+t/wo8Ud/f99agXQyfmppsEbrtJQY6KlYvaK9X5nBiwD+lKTD63kFCXX
mEI5GAdKZZMvIm0a+9gV/Bmt0pIPkNYVlllki8Q2iRWgKZp9FHz7cV+iy9WnrSdmLHGRH8/BeUE7
vnGplXYPBpH2PLqXWC6Z6RXmZWLp/O5QkhSJINTYDkEt8PxSvAPJVe5zKgiFvK7obh33dLm0vV6i
MLFLA9OhLzWbo31XtubsDHBjJ0+OM+PhD6oRyXalaY6Fy2ZcrFzNnQO5ASsXLw02Z1TX1TtzOOy7
l6yo/uXilLxmdUL1iwQ0DACAyWIZNig1WmAIXO3DkWTYUlCurx5PUeUGs2iLCqs3n/ZDyrzLEAir
wQnm2z6RDUkCX0NT77BHLT+wvoY36GWiWYSwl2wk/U4nhysVD8FjzM5JrpDP+7tRpBJZXVDHU7q3
dftkavehgsRlgn8Bf/ibY/VV1CmaJTGfli/3B0XsCvYwgjM51r8iVIErFJGyKT374s7qIQjp+Z97
Pn+Jbzizvn0fOj5s7qc4PWKwQ4eG4kJYTF1wVuVg9fyqFs7bsCBqO5VhsDJGiYwlzcZuWpNexCT/
BzMYdb6uAt2Zrt+GeIJ/huE8YvBgwDdUr3xlZ0Gdpke2VHVg71ISsJMyauJxwp3iFamWVlnCGktb
x/A17mbmdN7Gg9fBFQ/Uw2ruI8ZjZEbHF2xWmxBGpVXFYC7I9VQaNDNS/U2RlhtJgHrIBNOUVmZ7
XvJdo4lZx3f+Sx+OvRzLjvkLEiQ1vOGqIgPsU2pu9wvVk4dqtYM4rAUK0uOTiXvBcg4yUS/v5UMB
Zx/GyOxVmfig02hpVTQ73rrbVYPTSqWRF5IokqbgEc6JRu/LgdmtYuXZ/cXCuEH0TWFa7Grou3jP
oi4knFFBnG3MawEEI8x/PcWG3hkmJ06TSUAwx9535BdLHnbO9NqgrDLWsVoPQOKeR+bO3i/ATzoI
qryAIpyawBbRbYUocWfm+J7eGJw6o5gPnoSD91usVp8K592B9/5tg+9kRsxAfwiE08hvNI5tKpz6
kJg71p91EY1cn4qc9e4y5HDoxLoZBr4+xp8208l9+xDBEhREqK5aDPO/ntU6pVexPq8u+Bnrlw7E
Gs0p9ATX/UQqcn9XuF19IEwoDDpNnIOO668R/623hOWZyeGROCPkrN+kC6qPxkRqKjspF97fuVuB
M9cr4LHyffcR9Xuy7AEa+Eg9sIuHXtmgsCS4RIxC3RMPaq6aQ6yruy8R8OBMvriKk8A=
`pragma protect end_protected
