
module adc (
	clk_clk);	

	input		clk_clk;
endmodule
