// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Gc7t04DQJuxmOVrB28I1+bSveJeF8OvW0Uk1qMK4nwX6yAUkQkeNziU7EXfiIMR9Cl6f+PC9EwRt
Em0fbK2ZZLxGYeb1L0v+3bJGKPmHNHsJRayOVnzp9AqJlI/S9MuLuRFtWOXgHKnM4z82jLzI1AQl
9Glh//RIexjLCLADAT/qycteo/YCGPrcH8x00D8VEk44IgVV6yWblzC3JS/q1Xf63p/JsLulkaC/
m74rVbQCYHfq7SLrM9IRZ8nEWYvy7RC9xb1p/AQRACU+OleAIFm1EMicOxaxEH+vpabEwdt0G8hE
wUfoxbC5d83i+HVwN5ryTuZyaVXfL853UDgYxw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VnznI1OR0McW5FktFTW1ZS6X7+fZNCWAwYDW/DDDyibVmzOXUu9yyV3NboW939IUxOLI1NrMzY9C
qA6eaT1Go4OJOhG+TOICQusQR0AHC1EHUIlzbsjTMFvCs2/0+QASlKuSmMML9QHkVej1PWl/ns3u
kwjIpZkNBo6lrx/WO+qAX7UgiUHGw8jPYpVxThbO3r2PAyjk8W93SuW+aVYLMgLWr/Y2vk1E14/R
f6joVJAtBpSJ2/+fmdCrwVOUhTwmYPe1SN5+v7GJWwNAmhPiPSvxM36Ar/pEgo1BVvLS0tebRVXw
JL7Gu763JhTtApF5N3isq9zuEYuaFwMS7a3YHn1uLFCm9jnO4TdMuTjTWfFy9s3JMkskClBn97P+
YbRZItEMrWycMGc+TXAnG1itJePKlKe+jyZpluIzO4UMg7R+LKrIFbm1u9iQqjVlEARWNNrCqJTS
ea1GKj5h6WHFwcqo00Cx+X1J3JBejJC4ldnsp7XAXuTPqiwq4AHtMn58QNJ2dA3pHarbzIx0loHz
bfxFa8sOvOHCT/I6LhmLuhcMisq0PUafyXE53VYG3mrXOFJhAdNW7S7Mk+b07lJuMuGLUl4RWd02
QzZBrg3xI6zGsZ1PL0y9UV5OEFUELyH+QHyT1J6n7ODU1XteRxG0rLz/cIaYnTqxc58T9xvS0ntV
QOxoDCjOp+iU6PFVI1y9/qpyBogPS6V4OsYgzeVPtmvarGWRgDMHQ857GlbjjZ9mlboJG5bcntVh
ALV1QHtTtv5CrmbBd88+ofD5ldephUOu2H7ggDg0PBlETHJpCILjg+QUPZxqRQyCwk3lIAv19dEA
V6SusiV4jWsm/K96y54E09YHcB11o1Yw+lH4ovDiSoYth3R0A04DN0mYs1enyr4ilSKIuIJXWGB/
3z/jqwNr5efOSbHs3htE/lpZOwX+ebuSSHy3IXVF/f8HJfhgINRQ78pIouLAsPX8yRiIcObPJ20q
aT+0YA8OaBXTUzExf04kpgEeoUreGpVe7YQhtLQU7lb5zsvD4UM5RCB1SRII2yTjuRzaC2yiGxPr
Zxah2bCm/FlGA9IHEa3TZgtKK/vU4gG8P3KM/SDgqT9QawdeZqoWvD5NhPXoKcqpX92TePWS2HXC
/tsy6mvJAhtZ5XRZDgPLgMNJw6BJaSrlPNk+HcMpSWagrkub/bWYqKlLMzV9E5Fj4VrIKR1W/UHj
aiA06MjCASg9djc/Hh9NzZV+Dlj2VWCINSUwYHXwa+fAS1ajfNQ9MoJ5KzAbtLmCRNyFAxMGn1K4
RNTene8JKG968roDEDy435cmGrRbqp4T9HNlOTiiW8+tgvf+xr/GR12ztydI0kTBZurnciRvnCot
bQEbA4UMbn7poxRn5fLZquy62u/yQLP2kswQ0nfG03boI2yChxJmcyKqSXmbvkessuYXTTJVuJAy
sfFB5OWvHJ1IDK26l4MDTLKPqGZ/ia+++ji9v9jJieTf/ddn5RzIPAMyW16PQsFksw+9932g7eDO
HKqkRErXzAWi9aRdiZ48C1poxIAG83+Ok+W84pswRvJtT73sLK9GJQUwnUUgMMEY+Ag9i+srp+iH
u3u2mS046kOWLFbF36qNKGWInDGY0+pv/5lVPVNJ32+bb7wdJWYPt/yPHXG5FVPSsgHYVG8CnZ5z
B9qFbxyYgAHvTRmiyuZYw0A8nBuW44+h8vq8JnnimOK6m5jLoRkQuGVmdVLn9ma4UkQ+l9S1cJ6F
zpGOWSgCbaAwYAMGLc/w9vdNnkHMI3/K4CNdXYJNmVWM4/g8uk0yNrdc/iSQNQP8uxhbiG4Gg4S5
Q+spIWXSdJ5egC9BnJ5p6wq2fNsSWmvdCXVNY9MnqD7zYh5P8HWhKu/YjXLYAFupokD9Rg2HfgUd
DPw9AWevCfdjJz3wZSlhRO2h0SQd37aihI0aEfh2VN+drXUzjhgxeDSvblNswu0LJgkG5izPRjju
QRwXC31IA1qQXKryzWgADZLVKfkR1d0Qcsx/kz86uV4WYK+ZTS1qouOGFVVPqHUX5py0M8nLBcs4
nU3VQDXqxhbPn3gP9nrywzV4kMdHRILgnNApkxgYlIT2KOEB0JOmjDiEv7WN/nsu5u7Y8xHQmtr8
vSqNnZVt64Ljpss5N1yyTe8d46J0H8Fp/BvEIyi1P3t0LmLUS3iQtJm6JeU3YhB3BPhnCzn6s90r
5zBY8gkw0SHnUy1PT5a/Rcvdp8nUakMIz9ViNuash1/HKUv0ZuT9p+rYPZXb3gBYr8tkq8kXKcA6
TQu4HHtarBWnk14UTvvtfPpeyguSEX98jRt4sKcBw4ja4xe8XbmdJcWloHtSO4niZYJL92WxWM1Y
sYDzO6xyd8s2oMJpjNLfKI8av4uIYryZQXSM7llT9Y3N7Vc5xquMct+VfHaIVyah5Rv8Gj0tr++1
8bnIwpYWidMowdilkrbzQ7kTnYW5JxGm0GAhwRbkTiBkjlYgECaZm42qmdjLz5JN6alrUhVC2Ynj
pJWSxlwnfYJQMMfLOsMgYRV9GcBAhNSuPKCrhDmAcGQgmfmKkhtmKsxh80Dcmj4ticNU7uweXlNB
eQklocSoiO/Mow+phDb85Yj52UEqa+SCnv+f8b5EvfzOsMdsPmOz2OkYNsud3el5UpDrfWZznWAW
pQI0hqiTBwsFBhVjqD5tM8WjMOepaCAiKM8z301RK92D/T/l8W9Nbr4PvkbW5owyksaOs+qzzlSj
D5LTYkYQWfcl1Ue7YMDdTWzT8jhr4tHQWMTgE1LvdtsCsLBmv3lb8OzvXyId1kYmi/vAbzVjLqKu
n0oSGX2LRioG+/8TxhLrhm6vmaBmh0S6gGxX3S2BLFjYka5xJNfOoXcXU78UEUzAPN0HXVVFuYFy
mlpDFB93v0zGu2rP2cypSCOJ2g2wSbHNEOzR7KiLwxqd2uql6EwVRViQF/fEAx+zp9o2XOHf4dSi
N/3oSnW/ALtLyuyOt8aWGVvLfYKfbWZCjr/epBT8AQQY8TZRnYdMBguzAWtpubyWDSH1nj/PcoEf
UvE4B89P+x3YmpSVIaByEZxLZBqt+c8FZOGAVNgvRR8pLijYmUUCzW01ksOj4Cl8HKtHvoGXKiH5
lgDY16B1SwHHFvK2eTGr0H4BSkc5N5RZG7GAOv7sPa27mvqbLrHuEfMlQHNi6VuyqAoXKVvSmEC4
UHjveFK4UquENdZzOePwUuqtt7ugwVUkNYZLdp7bVoHNihMLw5aiTAeG5KCvqycUIqYkhDT8nh7l
avn6CAAK6pfEs8WqL3C3GSBlQv3xfs9FlEtZPI7zTMeokqan+5Ptf0IU7nCg756b2hPI+NKjTtGg
/wtyJCMvTQDFO2sPQlD1vJyPHx0rbEDlGY/sWpe/N6vc7pov3Jv89Jqnm+Q5Ptg4JFVP704Vusbf
6nghxgIfxLBfJzyVdW6CcZaJbExshp2oT3u4ufUJmKY/c2ovAwDLD1PW4awNWiqPYglNJuY4Fvbt
9kI7w6Hv/xIGaOnWGlkeA1K44Y4aXYHM5w1IYHNZgdrUA5+IpwtZP0DadO727S+roRzMTpagu5CR
tjFg+gMF2afDmuYIRxoFdydgPk9szG1OH29Lz5Yqqx64O9EmOj83maw23qOCd69W1jy2+UctCl/m
jo9qgXj+Uz9Oc2XSckQugsuGgx5kCsXBIlnef6lDfvX9OXsuUPeNHoz0M4LWjO1g0sXHTmMQuU7A
cUTOHqX3vrpvehR4q+XNJczbFGHBkRDOdDa9cnXsNg1QQhkGX/JscsYTjRtjzjtBBLRFHysS34tr
U4rCBmfGZSyi6G+QGb/xd0VFMSDHwBzoOj6IfIjx+v3VBDjZPs+CAwwbBKEJxVjxRbQkF7xXXm4t
kur32Nb2+Cl2aCyK8zSirjV4+4rXbK4aqVZKVezvBo4JScWs8jEzvUUbDLQ6u6yvWu2eHj6UX88V
yNXnqWwabEsII0PrvNqypMp3JQk23uYXlQp13laE/BSSHo5fJbztDK6io/Vtf23OV3kwaKAyiOgO
as6cAvSe0wshwdZXYZaDPq/FmxUfptooiBJ/utATj5EuxgkJpKx0mM5vJ+ki4w1lN7u3UbqVuooG
YNwY0C4+dOriZkZLeC9wOt/6UkDMfJdbPr2hUQCFoVL/gGBNQ8e5p+pLrv6g+38f3im92S9Y/4jj
8GtNsBUvcLGb7Lf7SVlUHBX+xLdfpCbEg8GIXyRkCZlsaZ1AsbxVMk6fl7SqouLa/jyiGx+RJkGt
s6zTxE7tHvwoR9XIq535/DRGLqjnSx20oRxRm8H41AMjjWR1Umf6tahlI/7A6vuDj7y1jaRq13hT
fZaxJyVCGsNiWzMBAnZjuXFsaUwtqM+uj3f8arSBqk6x/Vr2KTXG2/EAaV4LzrAzyMTtssyj+cfl
MSoUSdFZhXKj8a6MnpbZv9TKhu+cUIE/PZIQsRqzg41Wl4LBz6WKnoW61d/KvCKi6nTrdRu7kQHK
0ke9ofSxfAO4qElGtW3DV90R0/lFj83grEvCtN0NRd8l8zqjijZmscCLTQA4vkppoD/DRCd3Ob3m
5zRpt+5mECPfzlmvxYoxpOsltSaN6DCmmFT4SUiLXk+hh4+M+jf45RS9eOWtTvocBpO6to7uP9Ci
9kZRLZT70jOS9QSIhW2CZK2uQUHKdmUe8AI9wEPK8bg3FaxP4DMplD0coZeCCQS65NTBKz1RWCHb
IwHUHeo+ESHzZBAbVNCF6UUqREGOq9cI/JVzHaaRP31KC65pPi6U4twvJp4wZCs+nfQGGWBZHkZC
kgqS6Wa3ZVj3Wi+dwekfM7SQB79EzRJo5PUQ5dmClccKlLAYD54kiDX5rQn8L4FgcE1PvjK8uoN0
6rBLneQZC0taLEcTHhFuEtUHJJ7PjHEftL4//LyQ2QYTKzsw99WlP2ErH8tBq1I3Gxekz1ONsgRY
ZbyRcPXtvnm36nGzlMRzibiWGAg6c6OYnbO9Cbe051qKBrhcTCar+p29R4tnWgKKvxf7lW6N3OjX
bdhxt1JE+7kTtXyQ43bTTXJ4fqsiWCE5dOcRAY/VIIKBsN/dZO/0Av6fMuYyUnxzr19kiBksJbxg
iUVV/Oq7FWj8k0iMHyB5WSnKZv1J1yVkABC82fvPgFgoLpTxLdOW6QO+7XOglOGiOermEj3IapFw
llMIy8xdnpo7UVkEOnHHyym2LfRpkc9tRSpQ9sJHdFSGW5yOslrrFOclZ6N5G7qBcyWNHD3+iITq
J13vMXhccyFzNvEOJfEYjlveogVhvlCTtmbHu1JXS0HvbO0wFw3BYpp2UtOcxXbACGNKp2TZorL5
20B+T8XNMTMUvC+NLFwy5ydtN0deyjsdZjqLpoukzyYf35uYu+lyj8TX/7BC9BAxpTcOExFaLRAE
jxLwamk2s8zUH1hPgCyCkjbD/PIzgA75suf5yKfrn/1I5/64Kh7h73FnmwOPYdbJTT02F7XpgUhE
Lrp5pSCjIvR9C4sBundGWkM6EK/NrONhWRe3AJpqW9mtROhJhT5dJV3YReKG7HlpLfFapeyT3CN2
CnJYgSSmxc+Ary9tWZNAe1mP7uolrfTFx8aSXodC6Q9ugLe+L+h5pSNXI4n7b3AbAs9EubXA/d09
cao2+omh0lf3DVXMeMas8CUD8906tFSXiT3cpDJq1CTU096gvyKwev4ysv8eYxnL3mkO3UjsLVdG
BL8pfOopOp5Y4c5CkFtsW0E2x6y2zb0n1tlChz2h94yJgl2c8XR8stwubiqmKYQoaIFA3HOobL0y
Ys7HZGCG8+f+oc0uP0OQsj7OmnOY8Ac6oCbsb476oLUbaFsDm8Q2edVjoYJFu0B+3spTfQbLTUrf
2nfDpg7bD6x50NAaZe+bafPoyHBVfzLAu+HFKxwuOOAcNy4tQp8sjswV8N1cXvlvSdI1a21hfEtX
+h2XdGLDF0T9BIRiOnlPVaVh/jVI6cAvI59dHbUELF1FQbVoyqr17kAbXClCmweBGGXz6w3udk0b
jPuDr7MBoFGVwZ7T8nBRrAhm7SsSoR1o/d/ysmDaE0uA9JYgPX3KuBv6eyjU6xu9F9/7KIsnAG0S
gwSdedAIQI91cpDykeR9TctQRI1OoB2IPCHHRmt4mfaNzmpKxoukul1iuYfObwJ49lTXOAIjV2Uj
M3s8tB/5TBs8V7Z/DJ2AYqfS565Re3kEYrdmsDvCKV+RseMUv/52kW2obA1jI2dhgvg/zCKaSPWK
yJXYrmzeW2FU5pEYHudNP4RrSIzVnqDkRAyw6f37VGpevLk7qF7bTaRnJ18tgVHMx0mOWcfIcpq1
ccVn9ULQ3aCZPQ/sao0pu2Sbig3WhH8BhFs2D2hEw9bbMcK+9/HjguAjpFhxqMbMOJMRfVfKHngc
kykTXSS4RdnT2G/b7rJfzqnZZDR8q9tH0I6Fs4TndKaIyS1h5Qs+gWHnpMqVOrYl76loTyj5/e/1
gMC3cYcUJqEdbfO8vqYmiRdEUVwpdKnJD+C8uraSSbcrxwBd9wX3maA+vvz5WmCcO6wm0jNliTnX
cSq9oubkN32j11UIetiIdAZdcckxZRlMAdFRhOL3zGEu2cXGKBH6inUr4uZU8C503nnvpxO8n4vH
HPv/Cv+nz00cuMkhue2oBsTI0oFHmE+mPZuMv8+s7mO4BMYajhHrKw2Xcf1+9OMDnXm2wthaNfaQ
6e7gF5vHjfywEDMzXSWEuuUAD9/wdKi5zSTk9reRbRIzVP6b5bZUl4IDMzECx5kK2YAlzVqYUBiF
Twr0JQjaNxxTOk6YuaSBzUxrUU494vj98ViLfWrgzX46nBBWJYbYcGMDOQ7IvwL8rudB2erF73IL
uZdjassj/7O7wVXuUGOmMTeyHCr0Vz9gI+0r3ZE0H8odjqT0G1FKSBhQYLpX0g8GId0zifH1ZoB6
+6WQ/Wxcrphb+MQ1tI6vxF6znu/ERXpHHT5RETYQNXVelTAeB0scBDJVUlwOAeM6zXwn8ppPyBOR
WK7Xhgc0Ywp93YZETUEBY5t3BI95v5aLo4b2ufEDzOGJ6iQqWeUH7sXlkenQ2puWpN0y1FIouN9E
7vTMbJbBgAKeetC9z2PrAsb15orYTaGY2ks7Wc3mO58nJ3KoLbCuMA4DOVCDlzBBDd1fjWr56sKV
MSZGI/lvd6kY5XXGOmFXLmH60gPq2rCvQti6Xv+xsXPdi2ZlepKmdpPPh3vK2tcwpoPmKjiPowYn
+XmdG1dPrJHto1B/CThSDFIKyqdpe9u6rxYLs/B0EHDM4tjhrnWixgJOICnpLqF/nLBa4/3f0kV0
kss6V6kAG2VT+aettojQ0mtBU1FsSU4sItqqUP3TJPCTGUfqSxlVAd/+8NVrMzkjy6VJwD0E0Nsb
ZpY/psMECA6ikc1hYQ37C6L49PXS7yuoEVMD4VjGcwu7W/RnKQoGvBrahEZqN2v1T/dT5ClS0Tz5
AD0RvmVfNj55yWU2/qNNirf+6YWQ2o+BBWOFo8gR/6qhTeuVjte0GykICMLqN+Ef+HIJB30vx1zG
ACNyeyAbNPyiBH9Dmfz0FbIzEPqhiwi88Vve368vmCzocvfBEz8DH/mFf3tIG/1RmKhexYrHHi0/
NVcMQz3yB7TnaQALhcYaHoWxFDQiMyIeVIqHIroNGPBG6DJ5QEFwKkkkVqtD3XMjjKOZs0pz+Kks
XC8r/0/TkFJjrYnXPm17Q6UUatfcvGZFNl8njZ/U8ifzu5zKcjZ9Jm5YlnZzH6Arfq1dazF7u9Nf
mbwlnqIGYjSN7s5oIKqCy19ucbXyZ37oUvgEYbf2pYLUZp5YRzxWX6BepmFJm3agg5X3Hpu1oJud
ryTsoopGsI4qcBM81ICKQMcng5md3W/Cgrx9n5lrcIVe+Hwy1GsvHmIvUIU5FSXwRYT0Slk2WZfq
DOu8EmvZFzuRN7/YQJIMGZuXW5iGPx4F8Ae4FpW+SeifSgagM/rGAzg/nv6A4xC8kJMGIUBnMa08
4VQPcJS02hk1LXS746ucBSVB2Qb4f2QdfgsVidsUhEkE9BuPHN+syySqrVjQ7wRtqNdKDjrk29Dm
+l3PWTGjnaWHkrcKfG+OXI+ET7rrTlvXNOAOHLWrzOSy374Qen8wfI9op8Xas8OeeWsxZvc770cN
DxjyKoKI527tWsq1J6Z1fuo3/gkmEG37pN+62zlK4U/SboNSKFKUW/HaF675p8OLPB6S081yYrE8
rJK8wOlbkuTGSVm8rLXEoYZ9JxYNvd8CzgdrbaeB4mJ5/QbnBMM37oIuFDLys20xiPCR8Cosu2s2
EZ3F3VCdztWFNZXyasAOsEenq3qk8gj8ofbBgcUyIQdSY0qLVz0j++QHELuhwfHjaT/Hoxpg9IYU
ERCwVYemuwoRWtDTIJjJ/p3lBMyGAXjY1+ClAWVMA/SB12pjSkGwD7AT3uM/0EoeOXCH5vDo9ttN
V/4CPN2R3eZxerYrQHI5ib3d0KD/4wLO8nodue35iFGSq4UrrmD6GOVfU571TJ8qG4eXVKp6spCd
8bcplcrEgbfZ8PHiB+SKiJFi3mk9r9OlhgEJriJ4n0S6dLw04fHYaOcaIomn/bLDCcCdt8jC8i9R
xdThZ63PNods2rCrhr92sywGIxEE3VGk8CkpsO/ru+oIuoMzTDqXJEOhxefWiQvoEH0r1Ha5sp8L
NdJE0RCqaRYuWsYYY6L6e6H1B7IvBzxVgKjLLYl25tJmebzQbarjhhFbc1hb5PjxMgNrk91m0d6A
4rRbg43R2STL6x+Ud8jcIvElEPmwe3sKlLWCPAFVJ27cByeEzQAOu9xfEQlRTib7NjoXT5IdWjmn
U9MCvyeMB38S8woYLgZq8xSwJ3tySv9jJqdMjYbWKfmTNo+rPxIXsD4s6LK437eEZMnKAShj+Lyt
eS/MLxtJYAvHWlda4o5vKvKHA6r/IqtNlcLnGltkqZI9gesd3mCcEd5qHyW8BS6OGVW5vhr3twNn
KsAKm8aOiU3DyVzgoHi2NolrQFGRD8ylY36ubMVMWsWT4w17oc4CSxJjudF0gAFXdLoOIFP83ntr
4XpDGEiY2WaAcO7IoOrHxfDDxnUjWkXaPjyUsoAWrbFl2UXWSC91lItm2Q29JqjhoMwrm6RLrWtF
ZPZ0Fi+ilfcH7tOeT7ZwSOPxa4nDTS8BD6lZHQ7hpx2t9nlhNUceIhzGV8HGImh7VhCQUA0TnySt
I7++qsWYTzP3tSE+KM/J6y17aoXERO3drKnNKER1BveXeknGvgNtJ1ouDhmFDmmPc+koKlBOLf5a
ngwtWkDfO7wG7IECJco+nm/sido5DX+fIAdmNDL2g0A30vJPIgJDtnkuqytmJs48ZiUNMew7GJO9
q1QxhUQSrfaWZtYDsckhJ3CcvFIhCUKBqJwJlOEONNOnve9/nXpfCBBopYJYLn4VOXS2Arxs3J+A
ks+xuu8Zro53MJK/Q67Ka2UDMIK8OJ49ivkRsASWh7V1huigC1yrAMEg1+i76cCUSqGhaGRWA4Ui
rfJB42fWnpi0bSVz0kYyLZi6FXNBbn20Hkg/19y+TTA0yQ5zCnBjcKa6OkxgY4XGwNWnuwMVpCVP
rvzO5Sf3eq7+gAxjWzG++V5eL/7xr0dfjYXS7qnV7HyKiZXqYIYc9BGWxi+Vjv2atgNvhzUeAVUV
NUBiHsAg9Dhyc1zQj4UMvgqX653amqXcbRTb2C/36ULs+UAC+a88pAo4wgHfJElo/aJ5uSrvSc5x
apGRTriDEGgpF5OVmr9cUpvNByeEiM+hB/AZPq+f49925W2zdgZTF+EeFOeK8IWnKAFF7wjlPuU+
L0Ly8WiLIWHwUBxAm8MJhuxU98BjDInpnPWEDDIHYE71yLlia0EBKDRNXKEWhq2XOWbYOwvQFfRe
UHP1TYRDF6hw88ov97iIXANfeZ7Q6AVpxHyvh3Gk7qkhFrLEw93pem/8Lzff02+KdtnvvGNJmWhK
39puqzEgtplyGXTH7QNElTPbmgPQdQnarz5WRIofp7yJm2W5lkw13I4cQVUu/7IG5wtjsoSMhXHQ
ThfvhVour1f5uL3a81ckyTLTJL9+7Y37mQ+M6PSwpi12oOoir18gY3/HZZhyElF0wap5vRI0ry3t
4id1kh7ygeKGczuvCmKYewSoFAmwVAwvZSF1ViGq79XFkbIayXVZcysYlHVDX0jZt+45Fpa56Pvq
LIfbEjKJQ15KZLFyyE5Pvc1/N90f67d2vouuWHb+B6/jxtF9WNErHN9PpxxJRjy4/B8xxefqY/Yf
p4p6Y4XV/NltGkikI52UPRYF/t0BYoX+SATPoAG0+MMEGavJKjof+O1BvJxNthzIuzHwNrAwQ6jd
CR83lza4CAfWLRFOheKS7e9vaDbkp4i1hVlY0X9IuIz4IeAowc/bxvBTpUqxC0Gs7aTPLbMsVM7F
PYtep3wGHGWwxZGM9a9sPlGH5tWKM51QTjYYfcAn/tmsEoCxl+TfKubGm70GSIByZDkWMS0voL5d
dn7svc+kWzka8vOa1huvVRh8pZGWm+0dXrYQj8LOf64miWcmjvlBOunsBKjGPA34yWIIycoV8Hft
XzzVI6tSUCe5+5DT67YBnFO6Fk0bycskELd/s7cddfIomWvWH9yozaVgTVx999I3JF3n/hckoTD6
25+xsqTOA7AgmoUO6FSGEklYNyp1KK2QpXJbQ0MDuLSc6D1vJLa7EClwCvgkvz2ayjcOxFEmVWvv
HPq15WYdUk0dt3E+5xHFNWEmp1lKTio1T2SjfU/4nd04gJKRJ7HUaCP7Qnq2YRGuxdpX2qFWK9uJ
9dVFfs5Tg1IiOSHPenPMDGnWTomBmAlgjXCKmYUkmZ455cAPmIIZqhzqgKwsXIjeAmyiyz1X0LTm
IcUnQ3RUy6pKpKCOjzqkw//lDGiizo+ZC8Os0yqM7hDvOPb5I7uLaBm3iVP48sXj8Fu5lV4LhrHp
7Y9ODhdbu9kuyA8lian9FStBKYA+LkjLnkaWwmwLsEIZNLKenGl7z3UziIfLLRhQ1D4rPXEfNR2f
VbiuvsguYEjtJq4Kt/t2ouWFMADjyxuIT2sit/cnA3xUcr0IGQD1jtIdmp/rEwdLQELsX0X3k39w
aRU6TXVdem6lKzmlWyHF2BUCmHCH3hW4vPxmO4ug4TzuxIYqBkWB4BIaq4gQfmYEs8x479eNSQry
NxB7Ntd/HgqnXmaF2KfRdqLqWC0pBKhAbR/YeaI/q/PMClIn3McZEIPzKRvsgQdbouFkLaORCah0
/wqym23iNX/9KLnsxUf5W+MyEnLyHZcsBSuXRYVv4PpSXHw6T3noAQuziwhZuQDpJkJYf0EvW+2C
j5WXVUW6alqUxGYNknKOJQtRPDkZ5bMu/zbzNF2nMVdXayv0HP1YdLrJ2uxYmEJCjylX/PeyPXrS
py5JIJLt+/GPL4PRFuxlL+S3EX8FutdY2HEkFWoVWwjABtn2odsCXCksCcql3xjOyyiNF2qjHVsl
uCAO4KglBO1+22vRuFM5KQRvfRwsFm+TwTZd5OdAe7qA0/1RIbIPUDDQ8cXHyqbYLNNPpEHJXvgE
y/oJGOI0oYc30pu8bAu3UvOxwfo3YByxma72W+wMaeYOLcSnJTBj3f8AOyrBzcA9DeWCR4k4tug5
WEGftcTE3GpA4rU81D6zyofgjT3ZZ4QjeQ0EA9D8PT7Bs5JsPU3oT28J3bGPINgPHqe+uBvUgeRm
my1jd5mZ8SQUax0zZOB1ERy1I1XX0KLxMPMlcZoFmaW7dk0Y9enOTSzOQEZrhWVwjslb7oB0LEM8
knwhnDRpJ1mXZJgtPU/sVr1tgsH/ySO+W6DbgeCGtMxBYl9LIHb+6IIYJ29gq/c3PaPOyT00Ei2n
QnG8ndqVq2QiL0Nuqzwg/5O/LkxhK5kCieFk87JEV2YkO5kFX1UVbx1Gj8D3Oz1JWObOlphp/Oq0
IC2NxOKF3pQo2U7nhz5AsQgOO2pKUZe1xBwE5mxKkyUCAwTRG0wepV/MmDH44YXHFa43Q3eE1rpc
gANXmjyYuypE18nyTSd6pn++e4YKXrbqNiTyjP3+Ss2w+hPaolMu9kJTjDdwCbc8983e3Yjt19Uh
zGabuhuUqijMkVyUoCGwsn/GSjpImMmOy8d/CMsciKWn6VhaBlrJTGzVU/HWvN7XMw7dFSzWvWHD
L26kUKB9eNVPnJO/jt03TTQeZG4vNBda80DoTKJ0qPcu3mGcAhl2R4H4xk7JkpvSJuMA+eBCZB6M
NsgT6kAB0JOOfgfJ9fYB0jCISEzzRGtnsLxdflhop/OqgA/+VkTXXX0+t3ovWGQnBEMBweenpu6E
xhhcPo23B+F/nnDP3x3UKnQkv8eISu4LK4Q5LckAoNYucwAWAtGSwNfRzfd2rr6xw6jiJ8o0K8Zu
B53UbDYQLUbtl1pXkjEb5AK6NefU5VjSTPvELrZAOZxrj9tZXtfjmtn8Uw2EDuc3d7tlLXDudrc8
7A+VFnM9VY4VJC+z6mkln/uQmj+4YlFo1VGDjusyecXs/GqKdo9+1k9YemaAHukuzuo2oYd75m5+
hOGTKVlCP85jUy7cxIf3lSZ8bfukuWu9Nl6DwTMCx+uiGyQgUXVBzjbI8HPQQKRXD29l7T3LgoC3
uQnDObdSgxHghi0fWO8IRkQbWisT/iJweAniWUDbG8G4KfntFo+GiLLQ0UsKFMHjitlkeTfykhrK
yZ8ug0IPDQ2DlgDiaLdQ5EXIGv/6Hg4mUA/xuXqNJjxboWjCM8fqPK8Gp1MMBlaFuY1Os/2VDW2Z
nba3bG2izNSZEUi6FIzjrJvc69yaTXCtepJQ5xfvJsL+ZoZDW5uat9TrQSlmz9ntMeLVAa6AX9Zv
AUR4Dw8vwyCBhv6Bt/1t5grdTKp28yzgM/BckRW2KYRFnOF47gDwOoUc52meBdE7eP8RNN6b3SH8
RzQruEtTVGSwYs3+35PXG1fkVqsgK8NquuW9uwQgWXEov1/13cg/h1AkrQ9KK1KxkVwPFps81W76
/O/bQ9pGF86Vv/oTq+0cWLwDSuFDsyjBtBxGbzDfBxWr0+gvZE4n7gSNWiIHP+jKmo41/dtwvZUd
PS1THgiKO2w39BKyADJSn4dPP1lw9BFI8kEOzVqatBb8YnMcJ3ECfLehadDmafvrrSOCy9zJgVcg
6sofTduCQyN7W3Avuw0+LGTep9b0I48BJUJPWnzFkNY7q6xQzNVK2qTSFLe1RQazjE9AiqI78CUP
QZ21B1N2GTmueCGPjCKL+fVKrgYyGl6DBnMM3ZUhUOcEGg6ttXDly5pfsAttaURsWfcbs8U4JDI8
sfsbuWYHj/nA1AP7SLjkBlgJKW9fbN0Q4xFgY4Guhp7HLFkpbHrZtpfUH5TyotWECn+KijXJh+vc
gBInoKTRLWVb0JNyCeZ3TGjSJ6IINXMcK5++hFmjqj4qLWfGF/JLBuOQvKWk6jkW+AUK/dX7Uk9S
82kKY/NJY4vN+ciG7/dTlqXcR5hz0QagE8Z8Cn746O4GMrwO/aaV9/srucBsSjoOoJGubbu1zr/a
Rwp7RB0/CMG4eah250+jJyhXWS+3KD0BA1jH6frI2xPSNNnx2O48BztThc92h1HTQATf5jUY67wm
9lT7cSXxikKOaKwkhs7/obusOxVbrj7X1BZAn3CENObMXbVNSLpj0YgBYtw1J7A4LAa4XhI3D3n9
X/QkZFm/RHvkFXVYkpNW+OGB90v977yEdgGWdMOdqmCqJTDCCulLmdFboeH0ePPue3Pa9tB9Rki7
+3SzE45CM1f+Jy9L2z2BuZpTFvBRlxJPN5MOvy5Dw5rDVlbmulOIQK/IY2d6ydGi48Z5WMo0TxAG
u/TTniCZ6yPiwXClbB0fb8cHyvnh7oOi0PtqaH07UK97UBFr5IdJuapOEo6Wvk+aZUlpIEbBUDho
W7aUYQaTwmsAj1uDRDmqOSkpQFRra+lATBSTYEU+Cho9JkpilC0yXQpzg/l7ryGmuCne/XVFp+4i
dh86yfAN5fmkB94dxgadv6rPHhQVVMtWtyKoF8OeWo/fR8Vbb9pJgmE/+RwtOQ2AgcPuF8v8fcQw
hDStIWThAhnDxYkjbp4xaaZAFwewFeGM0ZqIaJ09s9x2iJ5IhtRdGJBQpeH6HRjWDFZNEniP2Yly
uhVT6JWdTSJ2O5+PmAQQbx0B2FoeNIfRJT4uzHZUmBhTagWyiQyefcFoy35GzNsltnxa0hLcM/q5
MIVzWLmVU5wA/VGol7j/hAt2hs/pMHfARM4ewR/gRqq3CJOsIK2PN4Mm3oM/xq7OrY3WNFF9i+pt
svBMxwaQ3i2HpuGOVZu2Yl5L2puf2aNNlRAd+BxdjpdxqVvK0XChFOLbd3Wed5cQIVomuhMIsIKV
zeIZpMVD9znEhAXW+F/rqoohL38e+G9od3e0OOjVNsvG99cagoUbV+EYt7Zhw0ffix8gJtc1dBwT
aZfDOaglKPfyOlBaNYLX5ro6+0dfk1LDpy6O1Kb26e5sWoSIl50COxTL5xXMI9atoXhypNWGeRgr
phYjooKxeSfDMjsgZkdpBKwQszcyFBH+WDAu8wTKWsHNOeKSpd4D4rXisCrMxOSJJ3C1Kped6Vtm
2UkNC92TUN9L8qdau9plPhSQcwHspjZBWQ04li64szMkzYrNUM2Ya4IJKqb2za5AdY85FP6AEGh/
Shm+TMn+oLGzx+i8j3bB9M0wIburxOR0szWyQgjnTE/xBvjLGTL9pvgk/CsvbDMwUhEzv9ZDuVXe
JFICKvSZyjyWZujE49QlTYeURBxdVbSaufxwVy5Gmo8ElMgZ1Tu0bthkefUERh+i48K4oDxSxMuN
WSOugIEZ7Dco0M+3dgXZ9pP4uSYoQ7iz42QG7OmtlNHS1//tibdIkNRxYlcJDdoWC2rKeSate3dw
YwuDWlY2v/hDHVIbh0xbhyXIGyaiV5Cc8wpJNpV6BKZUNSbgEi+Ettv63u6GI3ni8dcotJMGh/dQ
pGb4V+6FMFHu4rgaTV899ED/Yjsze3xEYs/L+s7YR77AFdrlmMNKWuPPrmGCWoXDsg+AZengX3o8
4znqO5ANQNTXorGg/vLxy/0Dl1OdEymtx2Aj/4XZbmncWEfhNG1F0yT9VXJHfWJk0WpDwFgrPOlg
tCJK2s9GCBATZW3dTvjaDL1Z/aiBNcBVDEI/Ek8B7l1ZTwT7db+m34GCooX5ShwIu+QSGDBh1bvb
Ykh3sSmCY2f262JZdQqUW+7SGUFGuKKTSOQ4sflHEnCQZk7vYTksE0hv71g+8YXtMU5AtaLB9LJV
F2zmiXlLx3FhCFnKCB5UpYH4kdNu+PxXxlHN1PAF143t3PW9aD3qSOS+tAq5jmGiOuf2Ze6NGdMo
pNH5oIp/Af1L7gwFV60uztrtRMGa9FrKBXlqMFbHGt0yl161bBY1vQBt34IQBap9QzGMRjSZTaUW
6JtNPKkAjU2ngjT8aFBVHjrqxUTy/JdLKNWPEExBaGVtzIyZVOEgDICYNrTGOTlVLMWcTyUro1+b
hrx1/HgNdgcdghugEw7hUwsIZTbbUFSDzYs0VgWVixwg7XJxWvRyaD92EXO2k3s2xRqqmTIkMUXs
FhLNQNILv+giuqw3RnVe2MBXSkJY+KMOXw0n++4MkMuVGdqsoR8qXVhoZ7WvWymaCiR8nViNztj4
rbG8BiCFX65wiSymU1Dz32pnu0aVXn/po9JSsbF5xiF30mB6S6gefK3Y2/ffwoB4AJyhLrWavv5C
cV7F/nIAJyngyUFtd84MZ24tLMejiw9+v105Jvm0S64mnnjj3hGrtfEUx+cg3bcjrEBsfbbt5vtc
15TrJ1jtOoq+6+Yfqz63o4luK2KRqy3XCbSKb4uwWiZICT3Ds50rA2zpeIcQT3BpLCz9HM/CZaoO
/yR8phCi9CNJBaQ1ph3WFu4fyKYR9Ubj4XPRYMfGwCmQx1wku1PXlcRY5y3vGqjtmMvJSk6C2jjw
zUmKLpQNw81kxFDAeyg01bpkWJ/3rO6RHr4A7Rw6erGLzhT/R+7s7jEKkTHviKqK6UEYlGXCWIk5
BAQ+rVJBjVUaIUvOAxCZXVci+Li2jg3zELfC3R6Oe8q8LURX/Ulh4BUbqXY4ri0arley2/YGzSuR
FECVC8lYr6R9SVaso/u0pTtDWjkfDW+040kCx6vB0VLpqafi8alrva5swa8NiEgdn7WukE2Dn+kp
DNvL2KZy+3UTKdbEJU1ZjcaSH+PM5f0Qo+HlMVPS3ZS6jXVLkI6B9fM0/ta7PMU7AipyQ8HqfNGE
nBmxYINym4IEj0xlDWTe2HhmLMNxZpqRNkdZQhITPUKSGS/R+km6e4NfV8E7E5/YE9nPR2gvnEAv
0OJGVPUHxREIxqZwFfbHLb6TSqJ56asp3yU2ckW6R8sBxRBkmlzsVYiI0wrb8nnEv63pZuU1XCwH
AguOFVgvboOR4AL1xT+bdFl7El8GHvaTAtmHCbT+hkHI91jJ9QrnengrV5dTccPkIegHN1WtULJy
RrGyLrT/q6I9FO8qjomiez5IJT2VKMVEkgGcN7kqvYCDDjyue3NLqBvKpipveMwh5tpQa1y89qy3
GhMiBupWHv/y0qhRUTYVcPdB4MBjE2D/gjY6zpHjgn4ZSvsE2Wgrm5jZtkdeESH0YHlfVVvZAlFW
jKPGSMOBANoJYC7LVN8o1PxMA8G3Cx8OMeBJDYVmFJvKD3nStUZxWvw0XrRCsEoB8UQKX2qpAjm+
Ih4GsPlC65i72j8+ku1w1QdZaF17AY1pKM33s3huUJwof5reeC5RK0p8SRppCiUCTUHCO0kw+97Q
UlJhRWi3WGXXhf0BDmgTxLLBMJGNWkQKidDiIHbFahbGaqJ/vGb0rEV+eCMZgKod/eDbzdR/GczX
FsXFwYzxcgO0hlye4AXbAxhWfWpYSR0EeaWHF3bR7wLKL+xalL4MHApkYuREL8fhte/TBP6DOEj2
zx4xYrDN+QftSBK7YwfCnpbWc1Yez7Ml9EISIdqjS06c/z0AsQFTwB2c5CPzyoeOLRWB6h+Lk7oQ
slFsW4o5nXKpDH5yEr67lS4Fkq8W/xUoYl7TwLh0AJmzmjKCMXqSakrXrRtwWx6HKWRF1jL0oDla
HvJiFMjqTmpGuX9bU+O0rURrComKlCSPtmOS9ghg5T01jeXZg9V2BwEY9OFkwJyERIZWFRhotVHx
VuKoE6/V0N+ca+iL4mQu6e08AUmQuJqUOmtKLEb/kLmPhgNLYC4sLrqg70znOS49GLWIzWBqccFY
R+KpHPsJplR9ZLY21kJy5svTLP+NVyPF+2oesPAdVWTYWtOnqnons2Sy6LDIFPTFUEeQ3dgcKlwa
bzZ7kWw8bCibQ2MRIH2hG+SdMCpD/VTW4LXnotKgPQ52T2XW0gaH8STeTe7kGqMZJbmx61Llg+Tq
Xef/j0StgSdy7MWto9klirtcje6sDOtke4XJKF2Z++IES5FQ7D+5ygUBM2bd7QlD20pYv8hFciMA
YYpCGi4kunaT561LnUuQy1f4oRkDI9hDWVrtpzU4TBAejeRwXvNPGuVSAdE7biHpdw9cShFRtYM5
hNLIpVw4f2eXbaOtIDTiIZtQuoDv+umyNKZHVC6P8L1S39Zw/4gAACpLjZXEWsDc8XsJiUQ0hj+a
Em8ZM11lEGBsP5HtaPaRNFVTjctknYKV1qNG1+N6CBtTaRHZhoiW5D7jITxNzWUdg9M9xWNPnlB4
PeJU+qLeLxEcEdk695rPzv6lgVI9fQB2FC7BF338H9kEISTZ20I86vT3RLZNcBXmznXu6E+ecAfW
9RveiZcuzfHMF2ICYH6qCGQz/ib0Q+xri0dUnOUoQX2gJQZymE5hhm0xvuDGOZmNOibt+sbyFOrF
ly83WLzKfptFFcrUgqAqXdxrbjT4zLlRS8gHhO7/H1zf7wwX0EP1ADtX4ashtuKY1/6zhndbqCTj
yhxPBk4lVTaDCm2acdBhLNEypW91lGwsORIHDoaYpQoKvoRFvxLdleoYSM8gwwbQC+ybQf3TXf35
Q7GCezxHrl7mgiavve/vbuaD0oXx8EgQWaGDyDqy7zR1SyaxqadgueZVnnV5Eb1xY1Fu7mojhDv+
rw8OW8dyQSqdsbyxEyEVWs9lDuoz5wYqFgILmw9ryspIQAJR6J2Y5BnuSvhfG4zc1lOjGPyBScnr
DcDh3UgE/FU5c3F7TDTMqVR9OK/OOSknyw1boCFcM864K96XG3qkVcWu5W458trrgXIU4jYk8OUu
FFqbuPts5CA784yCmUASRqVABmVn47YjFv9dRkJvR9lSU8fc0G90OBmiCtVPhQngKyVYYIdzOewY
uDcvoOEuVJBi1TVEENY4eEzRkSwBDrKhDYkmT5QcaGkaAev/wA6tQwniHEL2ImmKC/T2AQpwp+mq
mESB2TqrQay3vsQ8gnGXr/V8RptQMwZN2WiQvASZ7uTYqU3OeWRLXuJNfXjruHA0xyQunY2OSpk8
8aKh/V34Th1wZszcqKTVVIMHdjICRN7x/zV6xkYc4KibETjFn+Df1u84SFN06aiTylNzd/e0jkjy
nzDvbkw6BFenf79czoW4ZC+WGzQL9gf2yAeihgcjmLxA82zQCDo1LptkpM3Mgkd7MBuz1psAX8Hy
3e+8Q0gXHFNB57dDXEn3HepREe4sfUyFgn90CwywC/JdI0aOARYWwLN39WYy8HNqNESpDu0kPMQA
DIUdwu1UMyaJ5LlbjpmHKy/XfEeEDEn77/DzESEtJaTtvkQjhGhsdT2Wmsy8Ww4w1YWm4P70RnNK
q3Ghm0JMS05quku6+SLMB4HxGfDTJ4ST7h8slJve6DjV1NzCbdyFImfTC+zB8JqO5VRmo9lu2c9U
3gWGugZIE/WwIH6z+d+0y4XvdvR3/2pw8ytOd7STENHv/uQ+nINDv18IpoQDlHqcgVITK8Dwnnrz
q7u4Zdt3fd3g3CwmnFMMcahCn1kfAN/PSi4mQJtIZBT5jEJUsRXiG18tmy4auxMvk7NclGSgK0lB
0ESV+h6uw1x/Zge+YvR+Es26Z/dxdHzjl4o5i5jeZty8bt+EJt5tIUEcsejE53rG0AWhkxBy+VE+
N3up4G/WHgSdjpDm69wvRiAcI2fX2/n9KV4ljKmlGGdRatIzA2r7wa5+X3ZuqJYpdWau0D++qg0D
5pfFz9TdkoEFXrH+rlqlgYLmN6YAJeJtRngrDhct4TYg4/ij6Rf5CTEi6cthsXbPVr+HAcLf7bEZ
iaBBSIOxeDfNDbAS2BV3rGlpxx/HkKWkTBcifELwimMa3SvyK+WvcPz1dWUjM2rvsJWFUD40ihN3
L4xwVUBxIBBpK5O3WtvXhBKu8RI1bzcYUjiQxj7mU3+ZJKBBTwqubNryCVrUBYYDEmJ/WEaLeFby
vCvAoSErLin+nNgPaRcvKV/D0EIoi+1/M0UR4LaE5OK92gA5c36HOCLwzKkMsQR00V5X5hlvZpIV
7ByAJl8CzTInhIbweo1o7wDX78bIu0iCwyAVwlQGZ3EkpzpSO3cA9SV6ZkzmKO1/nn4Qs3boufUo
q8QdCQngt+UP9Qdoorqtk0WFum0kimkrrQ/zVeJd0mj2yo4Ef0cnXpxpiffexqsdvOOZ/C2MB0A2
pi8nl9CKKK5UHyiELUmCDZRV4BK/AoIU5puXciis4UIK2rZ39LtYqXcRpAdZjhYOTlibGlorsWXE
ML62JhqbNKLapFUpUTqb1GP7nXrdvt+C8iO/wJo7Ppl/jdvccfk5+/at6dem1NS7vSe8thGKDA2R
PH9nEGGesTpszcptJCLxdF9JkPNxw5wdnGqeuYi7zM1bVB4/yveJfmow+ey85PVm4tlubdx9ckX7
4RAYsN3/MJhjRbPdEfUq1LRV7LtYy48ioOwKNMvrkIYIMh9kO8JPilxkvvJBcY4lGY6tOOJ98xUJ
kzGsyQ3kEald6MjHG5OfaG4OsfbdJs1dNfMaKX3XUEuuylcjrvUW2qTBDpqkvTycS9dw4yucA/5m
htZf+ANzVFbG6a2UfsRgCcKQ7hlINNQevPM1GE7QcOUWR6QtQvxdNWaDoxND6q8v85y42GWImT6C
ceHRN0bB+LJfNKaTt46s4wmD5/FCiVVxeQ+RFl97/3WUvJIbl0sicavtNyyUi4UH5zRb1XzU4mKn
LjgHw/MfKbBxJhaaiwrv9Y7P82n9KhfbMRLBgtL5X58OxhmeeuVdZX0XUBWrn71bZtucqC/rfhu2
OsXkSn4kJJAySWtcD5d8jC2TWeKc9DtRbFlLJB8mBbL2Y5ClqBt0laQgYdMBs4vWuCpvUUsUQ4k8
9QpZ/d/ksLPZuj6KYoRitbn2ZV43e/T/F+iVeWKs164RE8aqtmi8q9VxONmnCHybrP546YGjvOtq
71MF76ABfu6cjwb09hKu3+TDPiv0EcBZy5S1zrUoR+p3HLJwxvpMPvan4/2qTIhqLdnZTrrt8oAx
w3nUCuIkpG92WOzZKns3E7DIX9KJgKq0vcZ74OeLvnpguC+3uxsWWhTVb+iWFHkioTscAxfgvf+6
DCnZh5Xrx+Gw4mWEDOfKmA6zdXt/BdqVteuV7DQ2K6A3McgnfgcDXCKzn/UdRfwv1CA2gQ7CIDHN
QU0d7z9tPdjra2E/zsyJN9FmMcXNZwZZC3fwOeiAMZioi3USsLCf+6wyIHhts0x5AZ59KrXDeB1Z
TIOlHP+KVqCehgsXAOOeL8GMnmhK2cjEn5c4XbMH48smUU9H3cW8DZiWF+KZpuw0luSy86rtOaVW
ticSRp3XLjAD7Feqk3HUK6qdRBDYwx5wlU1LMrUb0e0GwGWtwnE4xwHwp2Xyvps+hHKYoQUcUrbg
JXm+jQXDwcxaVuctYVTn/Gxk67w7hJZrngRwTNbqXWMWKUXqsYSe+UjXBcAoFushbxbFH9857HjD
WoI/XHxcdttMux1/YGwAiyB6LQBgBopIt3WtSw5L0jKF8g+dPkQlIdS0kChWV489AmotEu1fqHU+
5igq0XWf6il7YkbI131oeYNeFXSwjQ4bWiskzl5/2p3jweo2Xl4W1rmrO62I0pefCsqr8n2udZ0/
13A27XyGzk78uOy6jYF5vC8vw3xZmAhxF+VBgyw5hGEJGuniz2L3/UZzAHaFyZX6FtRx6x8odaDt
Z4+SOA06wnRPDChUrffHjYYnXI921/72xVUdrNAWpUHEXe1U58Nzwcx4O6JuxeTqyfRvFraDjOc8
FqZkiv0QFODuj8RnmTuwLAm/U4lDBZeHXE5t7S0cTpAparWmlsV6E+7RIL/K8HNRPxtdIIzMeclQ
MYLtWRXbPEcE4n5qNDC4HuNtxKs6ylqYefTtqC3OhoMsFzLgqxPjMw+3ISzkG8Gh3zEqLF3q4y/d
Ac+2Qn7LuTFD0ek1cSaPa1kc8dTGGWv8hMjylqJoYEOYNBLgQYhHXMEXizayXC4ofmm2g5ND2s+w
PdIzwx4ctpJ6fcDde/DF8Tzgt6HDx+xPDJ580ZCwpn6Y9KDElofa0DlvUwR/iV9XSCH/lXlsbfX/
HB1okT8uiwoTj7agD8VV868fX6gmjYApCvuQIJWWTuMKVgtkQiVcPxlDWY6a+mZLhxaJ8wpi6Wkv
VnptRr1GrjiyiyEODnglSjwPGsx/aRWLJmrexPSgLvTa7s3uLY30qf4YNBIO8k3vOz8y2ekQNwTm
j4f8DBpOU932my6XA3WnAQg0DpMqBMspsXo+0laPVJzT626R3N91p1x/659/a2DJ5qO0rq6zLFo0
OBdywZahSELHZqiWVw3vO71yWqcxMXjFOLZtElYwnlvmiObdlwmh8XgsTrI3uprdzU3lcTDUbJEe
eLh5ft/xVoRZDQ0JOD3mVDx2W7B3mAhcffxlbFF4Rl+UQq5okWbIMZiGT324hl09qqb6YFj+11AI
Cz3TITO46VAHmUKK10N5gNA+P+VFfSHBI7kfvuT5kSOZ/fQtyu2nT0r58ri+Da4DF76qsrdBz4XB
6+wAG4SGFJq+VN85OKmnDjgGNKgLjzM18ya0RLPpSSTWCUZXoP+5qApxhyZYQLapTz2mzv+Il+GR
UR5CEepC1oqqJBZ3rQ1Z9pb3D7RqZVOpB3KE8JcTx5pALJLAMQGeVXPIisGA9+xBMv/DJMGrvYbT
kq8glHhLkxVveuVOaNcfQfQYnnPyefHcTFXehEq6Km28jmpDLKwhokSL2M1qtP1Gvw6J19DSKFQ9
Ib4DjNI5w8CZAEbOUISGN2OhjWlRHqChLxjTOUVTCPQf7YmDfF3yzTOTf44qZ+RCDC4d5I/i88D/
k7dabwroffa2k5dR0hDI78epHvO34kOVmc6GGQ+yVwIlqIItSuGg2/ehpbPenL4RNBynFbU4MrBM
GHmot6UGhc6E4IqSbdYsf7bDhjkb3IuAv6go4GNtI/rzMIFVIRQqM3p+IUwM2S5LMQ2b+bJMC/lo
AquGAN4YMNccnkL0OIwEOUV2eEtgCQFtQJHYpc6CpENOzkAFhnduDQKX1pNvBGiu8Mmwc7Ofo5ig
H58gElCjtR+KRmg1VhGahjkpWTFTW92gdYL7gWloSk4ZCZR+8YqtnigotE1VacJ8OFb0O+GBS1en
k6F9XR3HHNxibKW0h21TyJQvzCp/EcGay50bo+Yc43mP4lTaMyMq0DfaAd1Ay5gnKwWC2kmfiQJ2
KqPMUcl2KIr9CpNBKJ5tphotEsZGDkB6qioigP/RAuR5hY3n7V8gDpAxsrKJJlAgj/1EPtNi3HUV
RXhtrEmGQnsTPQrgqpKmklh+b8Q6mH62B41tGBO8zHzSRuWOCvczD0K5zb5NypVXDmElLP5bbQh/
zPRhQEJmOrhslXXlifLMt8xnLz0oLM03C8Md0skAlDusdIo3eKguPhGyasTkaySDPKJSCldS8Biu
vuOJ9jSZW0XSbg/P87ja6x7nyU0QSK4z4ChNfvVrZRJN1o7nTRRLCrRMIuOA9Tms82tukDJvFm06
uxC/ZgNUkUtlt6lJC2HNKTogtBN+TBTGWKY7GmzrhH1CK6YYOQTESblj6YJU8g8MkleHhF7+ZPcD
qabaDLWgMP83lE1vZ6G+xng3AZJ3BlKJIdP8qfgWi98PfzjhDEk0quWDNVzvP1Yaoq+LfhW7jg7J
8T2Npxs6zKh+6VxotFjQ6QH2TgP7/g5d7GPtjW+Sjlx2rtTzrGC7BKtZaw7xiVfQJ7aadse/kWrP
Ji3pJZd72Akex4gR23U9ZCF845q6xXjEHZVKdUr+AfIHzRT9j/PqhmXN/xkkoxzxRdR2k5t2L6W4
BVCtu8qlTQNtDSuX+6sF1Z2clB9nGM1Is9HVhn9WxEnDQSLmNcsDVpgSxiESdPYrQbHiXP/SVnrw
YZbeCuUi58eH1cWzQFat4z8dYtRIyQLqsWKMdsZEyp2nON7L+lbjaj1+EkF2Pzh1JGPYV/J6fnwD
j1qiK+XwLM60kfSjE/trMNNOMiarQTbwT6MXD6rGomxEu9wzFljb7V3thCrCQn8lHmaYh7Dl8SvZ
UEU5UCtz91Rdq2kvH2m5nGhZKOndLJWCorVt5nhCRCVJfOcVfsvAibF+QS9sVuNxgFxfE7U44Y+Q
yY934S+H0EDvu0Z1UHCJheX71C5P3BG8Q1fGPWgId2/jqEjRWHfbqzMy5yETdKLPyFlpaIjIp862
U5rt6h0iABEpEesu6OdwubNieggvIuBs4djmWeMRbOHucPKF0bMcLduozTgldMgXX6pqI0LNEWog
lL/Mc1+wzxin+EGlqTuj8VfNci3E0CXV5rzPo19u74RFLq7KCkzxwJjM/xIqjKI7ZjGN1znUFY+g
k1lBghM5lOVGkIzBT1gGO7ZeQOwyZ23BkickBDuASuAzt3X9UyX4Xmbfex+pMlGt1HdhDF6Ngws/
xLehjK5Ssu25MmXdVSWXT002GTyypvyGepxhePtiGI1evrslmMb34ZPj5E/ZCILzwtkmNl3ROwhL
qRb2UOLGVrRV21iDGhzH9lZygLnzeJleot2mB3a2yvtBZDjHB89NZQXv9E8VjxvDsMgxGTI0F+61
PKuExcSZYM25xdj9f/SSYbqDTfJYwY1s0JNk3amyPGZXHPKgAW3KwzjKqer1zqX+RV+jtj/M5d2c
eJ3zo5Zgkycv8v4G1XcH2wslYWYPPwqXPQLuh4Yamo/QMi1W8MNlwkH+zydtBoMFDPb0g2jcNyWp
QYdPGnjSC1z6SGe2mZFDPCpYDdJ0GjhXAz4IHVEcYnF5K3irPsQnPx4nW22dr9FSHKxN6PxOAXzg
pxIVhGvaby9b71fxuY6MywTHkxelclGDIIyWIB/JmPV5IkGUzGPAS/9v9IKX2Fp85uRPpdlMEUpH
G0owNqsp1SCx6xHgZRfh2iUhkXZWw0/f3gwes2bql4zVRGjBdaQP8Tv2+ewjahh6TjaN4XLqqDlH
I3njMHHcQ3ygmM+eJplFWgV1C1+gnzELxHtmlR7a5kPyElL4ByzFCS4zbOkoMHRJpxqgbWyFpb9H
mwhy8/LRw6PQHUqbWycPBG6peE9m8G+CGotIkdlkWg3Lz++UfjBc8XzLd0b2FoGVCgLby5h5lyr/
7LOIM+omWk0OClGX1vd0pukDUGrPZyM/G8qhTIXx1uNG2UEdtUIFuPTwjvgXB/Fqvn8XIowe/d+f
gnqoBt+xRm+B8Tga069BJ7+QC/n6VVi6iEgUkSwfdExGuahHJqAKM8lIJ0y1A1KL4QBPwFTR5Mh7
jFattn9cwc02EihG8dUFKsCxUbn5o0yIMqzHdDN+sm9TLS33Zmc2aVLb5IJbvXmQ+rf4p+6VMR73
l4LOHrh2cI73KpoK64mZRwaDlIfBH1JPzxAbmwv/NJehrRg7wi+RSBr4xXqJ66NDPJnvVW7bxgfe
o5Nfe2vgsyyFEBA6a+jsBWJ6YluH56RE8md+p2Whi5EgNMTEvdOZnD5052/kTVCoYk0cIxmOaZ5C
bLo8cpltg63IMUUF+zSnbAV+Mm7l9suobDl6JGP9TRCFf9NxuJwegU+8TG5TF86vB2QOX7rBCRbK
YlzfvDG9WiTxlmlqMi/NqEhf54S3QgoO7Ypy0+Qlf6k9Pu8fZ8UNoEHjuQmW/hCP06rPUSBQFA7G
pLA5BKEtTg9CSNwWs8cnYhoTQ3mEk1LeUoHO69vwXqlThQUEacB0WH5JUqfL3A4a9izSJIedt9yJ
qfX9U7tfOZV5wbB3rhesbOV9A0VfUiZQ/3byPJP4FAelOyzUMo5FcXurxHOBEoQA9MidJH5HiGcT
HzzJtbUWk2EyK5zv9iwT7IA4F6GQNCZcPTglUseAyS99ittvub7KG3RdIUnuWuDSrtPRXDYyRjw8
1mZUUydThUZEp/37zzBDOO2o08L69JnvvqT1gyBgFVhsel+G6pNPh3OXb33y7ok9+dwf46KOYwLg
7pNThg/WIdYqbnvyttHMS4DNpAUAuX6E6NMsvm9znFOQNZ8n/DfOGmoyxRCH1Bfnwsqmo/GMrabG
9rjOeLVyhdwuqXGdDmFPgtHF3VYaaSisObA1ROpxxbO38CVV0o3ozyqC9CWpd3z5um4EG4w9JKEp
6S9xGCYxUQsS/RVZEIBCVuJtU1toXa+xjF/ZzGotCHt205HTzsInkap80wclCHM7nM9mOXl8Hhnr
+eMtwAHTVcy9TzQbyBPiYAUCRCyZXdrWktwCSSkLXpW0xZXlUYqHmK5q+4kqpYRM5YlBzLyhk5LI
yOOlOii8eO0fCr5BbnMqlLp+EvgwGCEf+uMUK5xnZz4SpsGOBYkSLcA6PY2+0g3CgdpXklAvIU/X
uRC/8zDAnEBXAiwsAjfPflv7Av7rE7T5L2otqaNpt2Mj7nmOdyIf/T2aM9fxEeFSP86/dNCUKuph
xYGZWIj6sBpyGFCXpkxnaFiHK0WDRxzK3+X6LBcMlx4FpqTYXuCm/ujdBrrhrUo0sB86UD3vzZio
sICW+pQqNPGIhWlMMPT3W3afDMb+2h1+KOgeE2SwopEUTdxg2F9X+aonTFQo6ulHiL2Y0+LcptwQ
MeFO1Vx2fhi3qIW5zXSk8JlDVStJrLaRKvBMQK11gDl4W1vRVT9ehcfCOW93YKNfHRjv/zMCmqhZ
aGTDNQwPd6HFDT8wu+p3zjn+1GpBUAoEo3noVFaoTD3e6mskjIcP+vdHw3htmir35MmLCBNETgZc
D6McwZQ5smg/tJpL6Rr5FRALcYAL48wYqDndeUhlvNlpVNSkRAC50rARMmW6p6tmT/mJIUjMOGhw
ofG3ZXQAb6qBQpzzf2HxjhXjPWWR07f4t62FKHbG5a+6UtMj44Diui1T5rsA8ZidU/o5srCb5tqo
aeQFKtZx7AQWrTqmcAzS+WgEXbb6a4hokDtKMLfBhhYcqpsssrRytnGwQY+tqWtPuok5UyLl+ydl
0nOv4M1RA4uuQyQjp58+os1fecEotMhdcaavyZ3JQuSDmLPL7ECwRxgj4bsfLiFFimCfL7ywVJVu
mKYAgD74er0YuGXU/oWgyPrj6KozVlTztETpF062x/yytNgKihNftTPk7ifPypgxXzbvwkBu3DWV
dyLfR2emqfKKo7wpu18hvRGSZ4ScdCgOkYPeq4FnERCSc6/qvj9bvFchcKjWVTgz3vO5VwX9HUEz
n1cmcBx4UIcYpLUhwRIM2slIWRpDDRY3bAOoBMSUcjDfxbkKckJfzNIwzhJ9YnorhB45P9Kel19z
XKwIa55nohWoKSwKAGMBksdHGzJxNaoyXxsVGcgo7mwM5xyaOgw41CtgxFJBSm4nzpuU8YDhsCYY
W7998XpCedoyA9fdGMXwalXDi0zAFHRXoCbTB1gEPSKp/BLzXvSFx9DsQDcmi94FxPF6dP1RL4sj
wFB6qFoS8lUGWzz3FTOSqWHXhzok4kMA+xB0Ab2z0R/2Z+QFtnQqPKXVoP9cqZf5VGaWTB2KtH9V
2oZGKgLib/K1ohJP8grUzjM1LL+8dBCv343lUiJqIh9VOW83Ddn6wcn93ojVcn5720fJpjeof0sy
FJUsbA2wB5N2FXiMRv8+GaB/ubzoDFuWd/qNHfbplDAfKfwCzrg4QDJL88IJjVJFW59wuXUCMCDR
IJbcHJyU2Bklp2JtF6lg8PxZQVdMQyMKY+FfB6J32o67AMKGVdNkkNVvHavSGEP0HwfkwqlM6tLh
IMw6X1KGCV701O0kvwsszAWhITnoMI9dJHlBabUTNp5EiqSoxbOwKHaKn5DPor0pyA6zES6cUVsq
iobX6O4A2CvC6GpBs2dZrKBPsqFxJFA2Si5UJgdkj2ns9Sw3hXSLuhIYJj0tQ/FsSQ5Tst2/wRJC
stX30UC6IsU/+nXNs9knHLpT0PoqUJ1m9WOCew1fmadL6Rf/6gPjC7H1envwwkg+qqW+ayxS9gIi
ean28IrvOCoC+5rJB+xnlgn3XLdpzV7w2AQWaAYqsQ1HZ/aK0Qms04xL32n4D5trW5kYNC+PIxaT
Tbsd/Sj9cjs0C8Gn5gOWUKl3lvWNUmdCTQ6EmUHyHE1WhSY8MTSkNEZ6+wVvqkBMzp3c5Q3gMLBT
t2YdH/Y3OAY4GgkzNt2Hkmlh8SegRq/C1VukXYafAJzl4aZYyyp4zhPYtRQnV5RnYb5lfspg0LIg
pQtHWS+1FFDHwV6Kcvhy80Xd0jXIWN7cWYXVGDPjKpLt+4zj6qHbbgkcpMNv73cdz4a2+iXBTKan
GWT5sE9amUug7LUUARytKvWW3TdVAjqK8gYc6wCdFzHx/3me6R1Z6SKbT3N2rksN5VFgvSg7mVBh
FCXwPBm1Wox8MatydH9vXQ4ZvPoZiYoHAM6nBxgW9beydMGtp7b/QbRV9IdCkUsi+dR9In0Tbd8g
UXIgNdvM5eY09/CMR6yC7V3PlwDHd4Bfs3gsnBxl51p9DiyheCAGKLcg6o1rnfLmztK1N5iNeILm
hqQO+Mn4Pdu3jKzpG+ebIlOv7NvAgvA5/ZNyQimgbhrNFTt+Tk7SrZc3X2V3VuU5dMdYPI29GuNl
bkCcoW5Ymc0q7mp62OymFDRz9SWZie4V/I3/cJcdFxyXc7AJclO9KkLDXG2+Wt9SIjZ7LIj8qRjK
fyUP25vOLIrm/zAmWZhkIoG7gC5iiv1TCuGXacBf+3QPibqtffQKjylyqPqUhKMTOjCSCjeN0lGY
GXjhMPu9FghwiViEexEhuzYUOWa21gV8fQ5jb5D+e7FpCsb/2ob+3Gh8XPuB7aYjdvd382zLLOsC
DuvgxSOD4jW5lHs7mpBLzZcsUz4KUvbWigI5RWyU0HnF8LaIhW7yN/XG8+MO4uB5cf5G0s+y7VIJ
mB6y5KU6spOJBc7jMgdvQbVlFl85ip1lRg8GvJJ3eiVRu8gArEhAEqvBUT++tUxidLlcAJKBynVG
/wZ1CNCWdS14xXEKm8Mmla2ig2nLoy6HzWtoyR86JoiE+61QFKVYrAIwh1Xp3GQNTcM+XX1oCWRw
m5lMmUteCuFpjrPY4HXY113l0uNTZfhn12U1G82pZFk70nja2N+VRPAu1kUuYd73w0091HBZWtsp
ZMW+oQN/V/zh1JAbOoO93mIBuEleCDSKhlCrd5NUx1A6YVB+8LQs/6IM50huUaxFjxmpYJ+n3+1F
oLor1ROcuN8HAWoU6WQkwkGBR4kY0c9dnVpUmu5S4/MeIxxjAUnh1H0PG2BluIFqhjOonLZ/kw2r
wnTWlVhkBwhMyJnCVyZz//vQ3e36yjaW3W9z+goUEeqRhO6Wj9RJH1ORarpq4ptIv40N/NQfEOBh
INYCb0HdmFImSI5CQ7pAAMUYlkfTod2eemqfUK36a9usE+RzNcA+Ny9/SnU3n3+Tr+V/rfVbAbDD
++vCoXY6nMf/4vn15ECS6YGLu4QGnrCUfEZr2t2QOHzD2QewSYd8rlC4kjdDBHqYpA9Nz8kZWuTH
fqLKi0WiySKHpW3dKVM8CrRAJKLwoBZqMJonaNSPwDr9+Vss4yg9K9SIo8ID3IRd/4dqyn2xZSWP
NfcU83+LsExqytWQQ7B/gOHT+kpxEmVAKAMExsvualXcd3Eew/Negr7zt+wYTR3HwAhKDU7Acprb
CGb4U4up8ehyLAcWJq94mEe9mLFjQEQvFEPaWNf3jwxnNAPQfW4mMHTtGNvKIDxsmwk/eihzrQoF
muRsedjUfGtS4KsGzYLlzjkRwnFHIbpfI+RVFmUoVonKdMi6Za4Nm56WSoNGJcc8mCgySRe4a3FQ
/Du53Z66R4fF+ht8ywLUV4YNSU4Og9dugFlrYHyt8cQuqwiXznJyNw0UhQ+w9hv+h9DwNdiZml3z
kXKxNczVam2zKwrlfaSbMAWutliu54p6QBpxi1+pVNYxIoANNN1+RuFxytoV7wKxPjpKTb8TKOUj
DPkDmltW4102MInIeSCuI7jdBWbKV0JAe6QNmtLX72AxV5DmgyJY67PnZv3SDWNAMIVGNsV/riDJ
iT/XxwFI29/mS2YQqdQfUpUCIzHd0oZaJfHZBhbPa/p3r7BBkmfeZgQe9SjfqPySYnLTngsdUKKW
GCsoq0XGcQ/UxascIP6x3qZ7SavYHryvfz10YTH4Y3tVro4UfOdIrAlpUw7w8DWt9E4OLOsuG9Fe
YbyQWODwsBFObieN8EB7DNfcEvRQqJFQY7ZKs9t1FZNbOrhNC2Pe/bxMOy2+0zULP3OqQw4tCD4P
K1gDtSUQZJYlb9ZCpz0A261XzdbxjXY1U7J9Y8FHQ080k/NomtmjmLz0qow4ZEmsop7jqwH2sgbr
aHh4eNLa3erREC5F77U8BIPnvO+tacuZliinCbNMm2D9Mc2F8idon9h2D0l0n4iMUIunpsQLiv8h
hEpQso3drXYA5DZd9hun19lsAAGl4J1k5ISTtjbDO6bswNB0IZLL2mFtNwhcXJ/RghozE9fCF7dK
ncDTQ8B8t0PSb36tWQEhPCwF0rHWk2IfGHLVTPe/gtsQvscEeP3e3fgzEiNZEI9Yi+/Kt9cQ1XL4
LJDddYpljtQfvPeDwvwW1ny4bllDMn0QBColFz9h8/UWNNB0OoBdWp4X6h78VIQuaDPvLamH95dO
iIEvxTcvjzDFLaiJjxig6h97zRltoUGVNaXBdF2cWMBjlM2o/0TVIMWJm84rGZ0cN85TQsysFE8M
4MrQKgmqpluFx9HJa12yfsnWIW8tFnOc+p/HPmuUUqUf1+Qy9YGEvWjNhaMQsJZyI6CCTTy2wZH4
LpyRAkAsq13feL9gap5JMJYfne481izFgM0gqfP2GLNqaGutuQTNNWSwfZYo4syhJjiZFB70uf+B
2/sEBwsSuJo9OFn1LOCI2y8oruY3bkI5OKRsIlq1JeAJUDNVVlPWTrijqJl5cLYVlHbQ/CA7rx0L
AVbq58nuw31S7SWelIxKH8V5OZ0AXOy5wVIWVwTe6ezmWJZekCfeF/hV+iUhtru56wNAa6/+5th+
HttJb0jAW4pEdfpkg31UwPg/jbcpbXeOFkGKI8mDs9HU3kKEuob77bjAjQWE97e/RJ34WFVHZz05
KPX+i4ERe2V72v20EZHrwmy1pT1z2mdLpDpaovpYUw2wEutKzUNZZ6fmpOWAIje2FTr5uIY/jmov
UK4gxPoidqwj+Rc6FevgDxKXOLjYOHvSS1Om1tSihceb3pKrpd98F75rM4zy+XcRvmYqpHmtAcPD
bDyRUWPAZKL6wXJk5FKlTJEQcbnrRHxube0RiVTpG9o7ZzUOyvXTEVhqi+w93pjmELRYhYCV4p8E
vzraSfd9TPTMCPwBtIZYiZz8fnNn9f+/l7qHUU7e6pNMzg2PkYbr8NDQocHh3gul2GFL+va45SJm
ptByr7tyhgHWGt+Z87TXjDH4f896bCOJYVUtr/e7TLP1HZdV7CdOwGM+1mMts0o6+SIz65+qNGaJ
PWuZ2uCreys+BwJPDQBvpfRfirnzUNvyOQRIC9uV8l2+fPwb7wbj4zS1oCqfycjHHt7YKPetKcQL
wwewLjvp9rJ3FrE1aj/wJ7mAnFv69UDZZAK9TGX2bnjT5F/loOBlpL4iIqh4XOuoypX+Q1LhnvpL
o7lrrhFQC/68GNUwjHcgKxuiWwDqoCUxV06eT4jYi6pX8vyjvJ2X6wWP0ybIGMo2adtpZRHLcdFK
debA6mgzheJEvp+/fxpIijRtx8C/bOMrUaXg/4qxgCxSBHxI9OZ8MEd6eY+3fWy8pkE9Mw/p2p27
yPZlg7NILasaF3hDy1Jo2O1nAP7FkLO6ZZwlC4cSslgMqM0IpLg1XJch7+UZ2bdIxdS0OUx+q8UN
7xEPDdI5uytnZfz3k8WcgBfgu4RuBu3MnRO/k6LasQSof+tVLmEjozoXGHaeKvdA2kdjWYrAwmdU
fAjvkV2R799ipqmKzZ8T408yjQpJtQONjiqKwu3sQyDHhqwR1kwpSl9xVBt3NWMYJ1a+vFw87/TD
lRA2Vf2JOb4sBH6AGFxumys9gmjY3Qvw8Wg/fxPovPKXghxNir37ca9LvjHcjEw2reEHOEVN1Non
bI4Z/2ozQ8QFWeqnMc9H6pdFwvmJ78hy3Si7GeeP/u5jV3941LOuwcN7m/a4sFYjUqaqxHm4Wx5/
nDv0LbGFBrZ/DlN8wm+z7eynKYaD3M0D6HUoyTVBu2JZu/e9JWHv80OROjhdaxgf+ScIqynGof1R
j8Qf4XYnTAmDj7Z9gcVaraQsdTEKFp9+urktP1E7eL6LN8x3z0W20U37q6dpT+u2UEGaOVDP9bVd
1SoRKCjel2nJe0vBVmB4C2TlaqWsoNzaRyvQteQirgcj+ZqANBtBdbfsZ2Xw3eVdtCU6te19YjXw
mpHnknN24gv9tUEuBQIiGUrQv01Vc9bUME2kRT70uKjPMr3JtvUobVjV/9SSwa4aPMu6t849Q8TQ
azb+hH1q07h/uCwoQp77rlrEM8kHCiNcwps51UahY4L10+Zl7CcL+A8c8s6QxjW2YRvJRt2LUP6J
tTcZWBVn/yFDY5srxI+eeN5j7WiyjYe/uJNM4GGiqmcj3OoxJRvzY/OlaixCpV6sX0zV+V3wsGCR
KH98z22L66YuwHn35+GxdlHaf0MaeKfvAM9V+TOtTv96Ni0XW93A1VQnIExom1rUISmR/NTc7Fe5
YgmvqIhIzNtjOOqiNZ8ZRA9whSiGGJXjY1tD3wuwokvEegRfMbvTclx886z2iqMvdjb6CpRbKOYS
xbHA2YykO+YKMqScJuBr9bpHwmopgyIVJUmL3tBfW7VG4yGfaQJQBgaycxRpUR5f2HEhWD0c0MEl
YotJnA6ALgvXQ5/OGm0XP6XVfd638aJn4hjXSwoZ61zdwFoYWZ0wlKNldpmzine/zHe+5IYP9rZA
rTVhrhgvvQehO9Netlr2TKf7jQtOQghQPpmn78jUBWD5B14lonsEz8w5BtupK0Lo/WNTTDOawtvz
Nxo42jHq26fDGknHPluqbsbDaXwD3AHCJwqJajb74kzIKItkyZWst4nd7/ISAJGZcEhO0mxwl4AL
KtFdF031Xmx5j/KOM4K0UlIAgSyIKQ8wma1veQRMdPZyNCXvRoqWpRQZreU84XBBNbfKX0YHcoUV
w7hB8EvQ7my3hYvwSULWaGQ8CKO03YXbHTdd7FnaI9ZO2fEulIBCDCUTrzqOFq+B+cP+sL+yVDcA
UmR7lHF5RoGqAMn9nt589NHl2mT4q5rFR24MLFxzHkkKeb23Hp1k1KMciGs5HCZcMWi1Qum/hyrv
AGF+IzdWQDORKVAm1atd2MIW1t9DQo4kTWLIeIhUQCTkLMvbB0zhuJaAQBUYDF+9m3CKI951d9h0
ocis3sOV3sTT+9HoQcXIJFzh4dEjUH6/CYbm+G7xySKy1bDt8mRW/VF/JtBVKYN1TBZmtE8oGNua
YgU4GH2sSn3COErY0Lk6fHn/Ibny/4BmNqDq7UG33cgfU2Jj9zP5qfRa33kjZRNk+DrQV18reSlC
jGIKXWwehbnX75uryoEk04fBZXFgrxQhs/M3Dy0pucYn4VQk5tNx6NdcKyH1UHR4kGcKqeibFx9c
XqnMhFpS2787ptHWhevC+/+rS6lRm7nljyR0YwxEzk4xDPhfd30ozBeByqFsHYx+5++3oNurLx1I
f9YMYNR299fcA+XBtxcSAaDXcKGM96OJoFHKkz6PumXRk+QFjpqgK0avR70WniXIf1lp+Rb3H4MS
Dmzs3wyU0uS4JSoagV3iEPuQ+XE8e55Wc2+bIZ/B7glFiUG4RcEKIq9YS9Y698IwG5xFrlYHc9vb
t8qArI13OYAFcvgD8vzDVmgFLpVp9DgLRHRWaU3xhfg/mazy0vDKseNWwn6k6v7lXOlni2X8ABnZ
KC4nq2hcUeLHr5UVtZScR9KEd9c3kvqxC5cd7PGaMPQUCPYoH/QoIqoe+HcvO7Naf4XN1JW41cXN
Xs74v1N4LerHxA12MYQpd0Z2ezK3j+8xMF4qfkznehqZKCRPXdzknpuBtl93eaaHCe3BFFW+bNoq
nSjeJZMNdRyogmDszIBS2LGE5EaFh9/WnBJpJgOOA22HICtjnDeNbfhc6TiH7I8Oygjve+d6/p1L
E9ZlWVfKZrBvtH/m7Uj5w03sVIlOUobix9+VbsciyCpV6hy9zzcSzQGmnXTNr+JoKbUY+63Nhpql
uccp6gq0RqI5/FDcvqmrY0KGHWnWgosUuV3B7vqJk6tH9cqc/8rIci99iEGiDhCTD53igp9MwSaE
pxaJKUqv9ctMOBqTAaAvxtlUxonngZMmztJmudS3NmgK5j2UnmzaZoCUQa7Pvc4BPoiGJQjjdMTt
oh0FEP8aR3ZksDvpejHLuS/FKxgQ1hlbzwWQM5TefQ162IW85mYniJkqalxWlhuAbSjqe1j4ML8+
4GxN1bm5gbQo3r91TFmacGsHfhC4hGiNx556/KtGo1+Qf2mgEHN27Xl98STyk0WMUk/V3tlz/fl/
SOw6wQDMYXFZZ8aBK/o1o9UIlnR2/iA7d79gJI2/YS4pcFq7ZiDqLMfkyoDNZTjKziHHNhCGwOmE
LNirxTBoDxhXqDE0mojNVZkp8ZMF1lQzBnVgOxKIoTk384CwkZmMgsgvtq3Jl8XQZzK8QbP7sbAT
763WGj1sysIVukqRWxvFuvxZr6zdpwRCGJ67sBLkiXA4cuHTLDVcuooxhPSRUCcpOfusX80mMcBo
lz2Dbq8DnuM8bXL9YuDQzNOrhpCk+nNwvNv6JdPW3kqd6BdoFvF3t/IDZ4cmIpzY/kpDRo5WDDjW
Mlub//4bYj7k5/TNJsvjr9FpxFteQXU/Nh+99/s9zioDpdZFUMpnH5JxWOg68AflGmtoNftLrTuk
AzYkIMxuOL+rH7wtkfWypggu3Zlu+fLeCeDAmSmKtRAiY9gUeGlVSSwxDg0PJevYJT/0qPjfcpgs
Ft0IyL2Pgtkfy6ptmLkzgF9KCrw9wcDHYFaNV9mS7xCKtrbIVP6FpMDlmsr443cRJUPf7ED2xUyN
rjopV7Yw1bLGMuW06OaNPOp7LOZ/7aX5ueIN6Xy1egZUM8OfgpHyCX6NYaceoxa2sqUOhhwJ69rv
1xbycmbqCgiqvmp6knAINB9diVl7GgYT5dkpZbRkJkeR9Z8muA5MP2NnB1MnF+aqV4zzsu6fe2Y1
q/vB1eoBqJpjSd8sMKia3JWbWxgKtt2+TS261EdfhtNaGEmPkFy7M1mVM3FUmgZ+fi/nbPuJHRKD
IVdczclQ6FKj4qm0a3RqqLxhORpR0jULG3m0RP7T/WcROWGn7HkXvL/xeeldtktxUfv9PQ8bBKI3
I6CYBqSjuSOjth27VvDVPhye5DKXaQhnU4ljES4+6rsoKNeBNhdfdJydn9SoxyKz5yerYZ4GfyQK
TVlRQqXVLz7y1Tcd4zBI6fHzFJ1a92Bcslg+dNdahbV66tssbpsGltFMQ1ST2+PuT9/vMsz+yAJ1
SLbE1OhwevgPrdNoNLw+Xiwg5td5VTiY43q0/Yjgrc00IpK9u+vKB+Ul4jfqppZEYKToI08+VcDJ
fycssFJQe+KIymQBqGmmU23NxsJ0xDIdcFnDv6ZPU9bc5dLx3p22HEYaaGrnHjgmBqnRZyvPJkoK
veqxMm1QPEXU7sZw9NC0NgeXS5zahRwpp4YlCK5SDvm+l2d1ScN8ET1/QxLC3tWkGXGvVKL35bmu
Il4K6X5dpSq+beLQnLR7R7O071dSXzj5KeN9T8dvRymRjRN9++UfAWC6P60Qzqmx+8zxPtmX7veA
pICZkP5CwT6h1c27uvnzPISidMipaKDm9tcW9tie84HFRQ7nTK/j1adRnw1tmF9A5c+kH0L3J71J
4YvChhP5RqIAX6oZMW6ep7IQmHAeUjxsC0LXawg6HUxWvDgxYU/Qg7owX5NLn+WBPx2S50wJrX4F
158cMUxtPKdB/U6iY+t9FnQUbsWlVCkaUOlDjA9wyW9JsNZpyaEPdesZ/yuFndPBbfL+pH99gdyV
MdAz41DC4K34cWUMd7HCel1B2K5IRATQZW7qSW+Ce73lvfFIw/nbUxbn1qH8dbLrfmydG9f+unnf
x9qV/edCwXGw8iGbvbhzP0MeeIg14uQ7uIs5En77SNTmVi3PxPZ81/xvP+9PDmAVLarZajbgx9wA
HUvoVBOiIIlV1xfGSJMuu5TmDKWKvgHC6IZaefGe+5fpNCHYzgVkwINV53S5pXxyrZGbEGtzRYLD
YAt1l60l4kF1mv5TTvyheY2e4E0w7DEv5+jQulQbO0eBUyDpiaeqaGoAwdJXLJlV2hxdhl2uuZlq
3TEBGBscmW6Txv67SaTLRh5JS3KPizvTV7bw3y0DZIJaMgN1T1mz4cDV7H4IQXIDwIQ8PW+8i5Oh
/gGlAHMAX6q8ZswDHRuu1lQePQz92cjlAD9if5i1BjHyYopEigKfRDQPumZ3X3+d0O4ZDrCDJR/H
Ob6zJnMfc37XlzeYUQ69jNdz9JDUHxgrGB8RSDoSNp2a52WMWjh+4yvox560I0bifCyDFWVDcnfb
ankuZxpi2mgFfp3P3dmVLxQK8v/hVN0sG+VR0A71R4wv5v0aB/RjIvfYw2N5HHJyr781QhVESdpa
vUK+VDRHOGrJx9C626CAGoyjcZ76LC6oWMJ50KX58JQH/1WICEa0TCRNk2frauLNt7rudGDr2Zho
EmUCtkEnrxJ2Xra5A3rM5R2fBJUqUkPeP6L+y67RVc7EDU0PiIEyw++q7hqBdncUMPYtN6z9GQfu
2HStFKFXzpja9TUluQUb7qNEFyNf8cEsVIN1qSCm4sI9cG1NnzV+tW0BaCsQIWibmmFe4TlTCJIf
QMfwG4UxkiJ2qR79USpd/rX5tU5oe5SP/UFekf9tuUp1FgHoTHS/bpUZc48hUfc786YXU8IZpwiZ
3fTOivRS42rHedULbQHZ9QxQpJS8X3j3Msi22zUeZ8j+oZUs32370aaAJpM5PSTX8SnJOmVQYbdM
htwYeuoX1aHx1ukSd32vPJDsf9T3XpPhlTRWt1rAcqvieI8+LQ3JlQO4y5UIpxefJoNTFgRT94VR
NYn90QAZ+SPGaRB0LIB+eFr0MHNHXU9zaX7nKlcVIh1e087Fpj0J7dJGiYZGsSrQBp6RqJ47HlCF
g/OEwyrfLljM3RzFWu+6qZ5FoAqCWOrzkFhv4k4vV8NDGhR2S8hv4aCDuqfg98lV6My7ecp3wkhg
6sDunoq4iQCQHtcHMR9T8/97Tg5lriEQ4lxuKR3jMMOYxrPWjbnwSM2SUR3VPsSfIRTBX9iwSiez
k2dokijRFEmImQOABfDm5cqJdmqQHKOjTRqqY70OYHKjR0CSrCm8nHhwA0HdojSszd/EWFUc18rV
Pvs92jBKWas+wCtYJyk1wQopiaSq+sOl5iU9gWToz2G04bjYgj+pJjqb5mTO5F4segBnTx0CnGhO
Bs/6m7e7Ri8RYosMpK4z8DcBXzBQxNbp+V/LGbOvUJzuY4ItGkzxcFlJBPWZXBNM5v8cvSbh3483
7bw9TeDkx0ZBQYXyJ2baS62mIfpKjFFgmXfUPytzx28IA6KdrWK9KZV86q1OnBhaLHn/ZZ3KLQ5A
5ObW+RxEUl4Zkmz3hB8KTykcWuhrfda0Zgc1/9TjYAAohA4pzMOKb3roTUL5a8qKUtnS71u8GWrZ
h2I9h0DYSIP2WVZllgQ7VwaM4nJ3xl/UAAquP4x5n+KCLMJJScFySsVCekp/9kykyHHfAaD/gK5Q
XIScwrA0PLTDuIa6nh9GihhB+W+lUZ0SFrmCq4SAv2kSb/dQ/XHloyRu18s1prYQL1rJZoRJL/K1
5kSX4yfThhOALcMj8efo/rA1AnlE5EjmQqVXio4u1XRpKSggJDNbos+yUqs9ktz/wKDAV63Vv+5S
I2mYtqVxKBZWv9Occ6SNIA86p5Qc80mgIZV3uQ/jU9WXOvCmftEE9WmqqM8H/uY8FkW87IOHAioI
HtKmthjprQBhf+g0MYVE2HZsaEVoxG9MRS3wJpr8vTm0cxQGYnvHAMguRSgHUDNjLoi0dFExj+p8
08GWzY53lpOrtfnnARmaQfY3ukt6K7zFeGPd36jt9RcobCrVzBQ9Zebnpe4f88g9upiZ7MAWXUL1
JRsXGxNTHtz5is13rnjekdGG8ZCxbRmf+NmVr7leN0XRKwBzrtRdzdDT+h57mSEvuxYUaXd1B9gF
xXmmpPI074ofZEV3ugOJA4TfSXPzNUh+rO5MyOcv7CzKrgaqQzGeuiI+R19ssdCK3f3FZ1vT2unY
1a5xR4W+TOH/+W5BBBBlD8STptdlDbfYRgCHzZIDYjWD1j09AOb3DclT22jlSOz8KxGpjedP3vY0
WjXfgHXhcPT+JfeId5FuCNzxbQaU1qLA9KO/XZN1NH8J7u0wg/1Ja4jafoRn1EYXOonwts/5gkzT
WdcVVqPIRdnmW0gxliU0Tae+pCyEWFxun88BFD2qWjtvoDhZcW6LKvaA3pUfsoUYVUtcSBFmZygM
IR0+PRsIyb/evcdR9OW+NXJnTp5s/O+BZeuaeQuj4kq4+zYhSy9N6jV3ghQ+rpYkw/iWdFZvyC02
nIe+wg8Ct10zcUA9yrN/bnZRI2dBELWIGLI3C2xDHjP0k4N4McBkCf6gl5BA+nysjouLVy5zjrV4
WiPsIKEgGeSzV0oEkNYOZ6mMXrp95/9lr2Zbp1QjWAlWujmMOPfH0OOR8ycTo6T68LtT44EeaZR2
dVK2np6/xUkpy+gDbCY+eZMaSOKKwnKOUwahWl6toAvbkWp+Oa2ckQOHpkLv6q/EiWw/+YzhIUrH
V1HI8vYEkXFw3kl01WzWSpmsdczqrRiBb+RChZ3v/oqZ7sp9AiCsYBhQvMBq1LvOgZF0pvZ7Lx98
12WfPv5kV532hGUwUSZBUAHwPeu905wBYVOoNlnfE+fvLEL70Dr5TPw0zf59owC/r3IeXGdQvuem
h00Wadn5KWtTfuE6dKr3UuS1KTaHO/meX4GAW/8pX5PX66oQv3/HLvKDmhXHERTPsdBOqm7vicu1
W8pTAnx47W6B/qd98r68rsl3Jc/0FeBSvdX08Xbocr8OoeDwmtHIq+9+p+Cs+xHYf/M7rA5Yb1HS
Qz2Zi8ByY4l7tLp/AH1xqoqOAWovOTxcploOdKtSHv7sizJuQ66AKWPgZmhb5rjATv64Xc69rd52
5wDosbXVa78xQkN2+ftyLp23pixEZv3mMB/lH9O3MUsaIEKzL4C+Y1C29LC681u4F2RJn1HL2+d0
4AD2I+dIiGWoWI12YzMFGeUtcZtutpUBfR2ogjrJWLI85AHn43VQvkr/ISjtY7YdEtDNI0RthbF/
h7/hU+VirM2qeJwdy2FYdo9+F54L/PhxwGsEFTYiZJ92XTGQQaLqwxyt3sLl0dRcXV6Pa38XUMuR
ugc7lkLnbk1vKN4LLjqc/p2qkx3Nh4QGxLzsw+Vb2dwfMlujRGBiC+uyfo9nRu6Vbfgz4SvTXHXl
C1P20zmeUnrOv/6UsbP/24Bp/6zi1qco6rbpQ2lAsorKtiFoJ9IWwTNVHiYJp43wGyrcUxhPssCN
QLbX1/sAsh2uaulrpxMV25gyE82JbF3bUlkWq9vv23GOjrCI/4VBxuLcgPR+ArmODMq90pKSJ3GF
8vDVg0AbU0RtI20g/0z3gySZTKxerQ5ejvoDni5Uyqm9BYCNMP+ZsUKdKZdGDDK/iLRIUlKhW685
8tF2Gc2KMMzoybqDsGqhu4d0/M+bXXWMyerYz0+UZC74PZ4cwKFI6b8SIeLYWF91AbnH9TTfoa5N
byb4lX8G1L6bIvPNq2Jvm0FHWr5zf1dOkh6yFBPHI2Ag/qEOxeNY2AD7AZLn9GiHEtUYmfGJcH6y
c0xFcLrrW3YHyiw5CtdNfPeH9kEa8+NH9dQJ2b8Whm6dYz1paGVJztYcs+842uYSr9aJ6lGEN0+0
QS5RgC2WucXbESQO9oZ9BJxh5oUi0Rs6g9XdALEn76YbJS873ExteRqt50eYqz5b9xGQU1AA51R1
CT7OkVS1fgy4MkFUhn1WTH9TAsTRBRRyROmtd5S21pFkXGXY78mCG1kaKsiCNqclENTv581Mbxb/
061CJoY3dWyONd72Wyncg8l7AIunF6pNIfIM8fChOfyRl04zHyuE2GvZa7o2OaBLYZr9Q8F+JZRy
3S6cUFnyNSYTyljdXRhh6dvZA0wBt4mB4S/IYEbrgixdMdl/5guMy3AlCXpf94WQX+ULRE6I/sKP
opigkpauhhGxrePHnC8VLXRjCvMsPhxQx1YMN/LEb4pOTpd755Vai7u/GMFqIRuSOGerdxlmTaST
XXNA4NOFK1+kpr9dyZK83NnZt/zhj3Vufyi/3FXzfUEJL1dtJJe4T/dhFx1A4j6sXHdr4YKXoU6N
uAZ8rMksAvMD+xsWuHTtpw3OzckGBNfsNyeisyGivYknx52fM1P6CVv8urnh1BXClouxc6UQhBqH
XhmLN22sJsRNH36D/xxsQDy1RDXOeNqzf++aEhJxQykiN7iTqvSRX08SAHVFTRQwjH0xUOPZNQ5p
kYtlJSmn2u7hevXv7OdDBlliiVMZG153vshJrJ5KWb1WrASQywHVtdqeK1yod0SELyu4NRQlt8uz
QHkSTPjFxQMQX0zxU7Hc1RggMW2vm0ZZ75R6LbLyM1JHjl9OTvHmXmF3BNzPZuPu9SEjPAGeVzO+
VCYWo5EeIEvkK/UgwBE8DHRzutNWmD1FHu1O2+JLkeTqUOus1dI3KQAEQ27nOsm6lvIoHzFfYDPk
DjMSknsBKr2XPL0RITYvJOLrl/BxGDGelbn8NscbWEBY3ZzW3pWW8VxIilKFu9Vs0O7NkiybHl+b
quA6pAJYY0f2Y+S+vkou8hV36MmDTYDHqqB0Q+8dhMDQJVUCQ9IGjnSJLaK5wjSSOX0lSql7nEQu
Nl8x/QlOBAkglHBuQF2gzDANWpceU0AkvXf8rcqsgBnXdbXkRm9gCBvHcStRboaLNIT0BiswfEQL
d/pfaPFc1r2Eiudp2gK8eQ2qsFl30+j/KZ0Ui2Gl3oBKIP+RZ6rysb/z7+xpNYotoZH/WG+Bz+h8
zsh7tYiCm5EvDBo+ZYzvyXvvg4DdcunImf6LjS6Fomgto4Y7yo/RfAVB9akpn9dlJy7ltwDVjpyF
kx8+An8X6NCoI5j/co24B2ewJXOmWyfeeLH68JqBvPLCi6XeRrsUua5yuMagYrnefT59lGBUb31X
dh2TkFg7r/EJxdaK48VncyY5s2DBNMThCkTFryQT7uFkHBW2wFkoD8TWEe/OT2Qn5eXNWBejRMCE
dgY8feH9LOEM2JvrALE90TfOY4zoyc5o1sIKlBp9D0WWf9rOHbdcoS4p2ZuyV2N0StNZdkgFjyNl
NWKV+LecNsWz8mdybSVYIz/3N4kKk/kZVpEDtXDxtRsjwnZyeLF1Mi2PZxhjjKQ/21p18ot6pPI3
CWddgAUmKdKvzlZf+fbgx3BRmSRp8QgDZLp/HqhHe4aBzqh6f16VUMdtWsDnEbsFLFDZYvqqfCn1
huQLxMiGo6XyqdQLSw6j8pgsAk/jPS/sXdFSG/UzStz8bB1HQlA5+FwMmvhjmY64A3zkvXJRMu1b
6bkXLae1SUL7Dwv7e9EwxZbEqKPnAc9R9p+2GxNilGFH9w1LV0XxuizqIuiR1s7tdwUQF1JQw/i3
D/gWquTsQKHGyijjSIS4Ay/B6EmwL5iveyCmIap348i0qc5V6e8dhJZvTjGDnIhX4AdHyeVMeWna
2tWeELASpqMuidlwhkwsHGBxKLw7qQe4AcLWWS4IX/QRSv74yzPNvpgTDQ9rcdBXmEyggiNTve/7
QyP6AsJfIu2ATzx7ZM7LfSeJJU0HNxNt6JaTEaVm+fQVYT5wGMs8MNpTw1xlYCPWTevzc5wvGe8i
ZH/lZ99M2kmCdMy2knU9Nn+0IEBT36dfxOeWOOH1eFcVHiuesKVosPba+0rfVulGbL0qOaQ4yjFR
T98/aOo34twuF+GAW9IK57TcZ7Ejx00ccJQIlOcgoYWL/MDrRRJaACM7D8VW8QyuabOHbqRsj+ZD
62I6vR2kpApky5dQDA1nHEQui3LyeT2T2z5pqjAk0xlPQRR/abZSoRr0iUq2ECQTPSDG+6+a3IeJ
eD4BbiEJ+WzSEoM8j9P3AQkMLs0qK+nAHyIWobCffVw+wQYNR4RtiTOOBZTGB+KMAEDuEMZiYrvO
K8XDwVDBq19eWwxREBWYV68x34sKY6iMXRzxpiXsXjA0F/2GPki9A503q9OoEd74S+b46vDvNMVa
FHQEiWm5TDJZi/p2CjqhZJ5GZV31LmdYsl+JUD5t7K0vb7YOrlL9Jm9o5FMZyDJQ5aS9/4pQOP4Y
EByihXBHzJiyd7cFUSTftalrA+hubjOmlfYW3FUhLaWejnKYfpF+ttQoYkbs6oY6Ow/01nm3P1OK
oIZQLoL7OD1mHhA9eChU7X6EWAtoywNtDMYSJm+Rtje1pBzAVpV2l9Z39zqLb6mYMQcAU2Xe5bnx
RURg/IOxDQ5wlzRdLGI/9a7w/J6cKF2jVD2KW7EoQoAZm141yVzHCs3S1R8D8t82NMfhNxYDsw6T
03zf5GvxQtdiwMgQ0LdSw6tiMc5pKYMkRTpCv/NP3A16zyFm2j9jJo+wP1LlzlrLXPwFlCyCqbLq
G1VLhh+dFd/hixDfqR4QXVtfSODDwvCFhhVKpbb9tu0qccECkBBA2ne84V9dRsA+JtZimUAQ91Ei
iBBi0IDTvlkiURWK4+nPWaiNZxPFoAv5lB3JSpLUDFk+OthdZEHwsMN55hbf4uylB4J/Hdhw1WgO
eRjCfa6tf/qsXfQaKcQy6v6PwNmvcdWWSisUnebC6Uyi5qsMHYs1UD8gSt5yNozDqkhIxghHJ3cP
cNvC7a636AuYpGK/mYDLs4qOGjFz5FVCrp+XpuAwZzbvWhQEFH8q37/26GObffjvIEMMWrKiOvIn
wJqNKBzukdcsHvbrYYPB/I6/H23pPA0IP0GMIwMEu6pPtiers73v26b4NKL+Lmw8smLnSUDyWn1f
ZC4dMosz0FCJDrrQtN4qSOVgZ7LRMY4lLWRMi/ePduWxRV6vAhKGVjtpLcsQUDv8cM3ClShEAR14
+HRZkplMn0lE2fEmqWOBpfU+zmIksJzA9sT+dMmZNhQmDM1e42WweXgtEkOzVm0NlRI7ypCYHQpR
WOUwH+hMjvQ1dsk9rTEcs9Ge95sN0ZU8EWYIz/OC2BwhdIcuh1y/QrIRuDm48MPQSz/gSAquWeQM
I11w7ilywhgM7af05ukNThNBC81pkw0ku8YTY7IK9IICcs+L07/F/UJsk6YNNqdnD4C/D3LeAcbP
pPrveLJfu64NDNN4obQDcS2rqikeOIWVBog+8BjugnY0l5LIYVpo5H6EJmkER42qczcxkBqU2xYn
JMXF5NGlAzXa4t1nn/itEaGJkdfGQxmg/0DE4vFUMrDHLN3BBBqCQ/8Im4VqW4tK0KvSg6fCbjeq
zGNdYe3tdC8w3/yv33ThedCzwyhQy/PrnuubABbw6pTr+XxA21pM3S1q8nnnkrmA/huX9SIW1Pnf
2zHAan9NZEZ0wLU4fD97m8Suw6gnERJAmhdpC04LgkNjNYieKtVQoG/CjfhnxB3X2vZPkFaRyzRZ
dSdQIMspFGb47E4ZMZIFWJL0R+EwEdZtvGTqb1E8l5LCGT7xpqkZ9PNcBbIdlqzyJ//WPp8F8czR
jiz3FD+c+HbV0c3tV+6y/GNu1L4K3C0uBJLqyHG9zLoW9T+EOtTmbvmTyuWpj1VV/vGD/BjvYrou
IhXw6UVwVF8fYUdUSqDkGOtSHIczZ7bBD9gIyMtVon6aDIAelkOxflMhlOsE8gOUt/ZsFM3mTDIW
3HR+3Vg4ZH3DuVp6q5GLdIYCFj6OrNcCHuK35WejyYg9Ie6l7MJbndGkRhPWrzgdDHrAxWImjGDG
1wRuu2KY+jl4N88otUrE/GxecdxY6s8sWAsJoQ+kkbu0hKC79Q7D5+ZiX3h4S6za3OjnwdT7bq1C
ZZkFFt0wBVQ8g1kg79UxrSlg9gYVDO2Zml6xYrhAVNst8xBOvLj/t9pAaRX54jPHckqPVq9g4wmM
PLlFfayAHa8XGn8rN+mv8yNDfedJv+GyAlc/vaQvmNZ4yJwAkciMAxZVag8mIZcTN7iMa9ZKbJob
7eiIgOkDMzRPPKd232GkOgUThhLz9P5z74Oe6ELfbY/+5ZO4D9Q/+dbReFtftJSnoUfM29+02/ZR
IJ0Ox7uSrU1HelBzirW6iOvIZeDZaAHwarzLLVnFsDLU4/Pmvu0CniILyBqgNn2dF9qGdnQCYtof
KCx/TOARXDVqDDX7fbE0fYLZv1NoJyFQNM2v2w8vb+MZN42D6oUUlKx4f0yrqT4IsaGOjXlFe6Rr
ZxoVVGehwIff7k3hmaVDRKzNAs4hML68NBhSyxZDRyRIuPTkgaM8ttRgfYCvvzPhC7gDkzapzNvD
HR7luvdN4mSxAgxysdU2K/MI7D49Tn02mxQ4Fnmc5EGcq/6T/BWBMkm0eg/g6aQOMX2xNj0QxHww
Jzb+R2DUN3jPMYLF4eHMmn3eeAyIjbnzjJq2YGQhoKnElu9VRhziyDtjnS+hUNOoq29+HfWzG0bl
YEL7MvVTcj5k3sQ9CMlCNaU7vKE8zvBGgfeQJzdg3myEG0onHiJPDzj3RrMFr91fNBVTP5ERuoeq
IQIxELDcj3WckMZ7vjPQoWuxsi3Dl/xbxj55MPvzPSquLwSY2g5meXYO1xzZv0jc2exy3c+eI9Af
RI/BmZevz5I3DHDGUc8b4fx11WwLws+Jxpby2Bi7j/jkAEv7td/eX5JwPjRbVyOGc+grkiovJKfj
1yCv8qo43dt4AdnxjlfOKySj33sTrdTpgzNQzamV9Lx7ZjjHcQ57Y92TsBoG9mWYRl7ux8NjTHyw
jt0xUCMXgHaoyT4OAys39ND+wWgFFJOFyDV5S7D03wGf2AXp+SZ3LwhkQJcDXVpsTbqfM3W0w0QW
WZDbx97QruI+56FJpVoOJU4cTG513jo2rQvcYGf3cFh3STv/QyvbDZjMFcKOevQOXZKPEjmXVSrH
zHZ4YiA/80ar0HwovRZ17MjlZxdt63oIdWZHvK5rcJgdwFN7wloEq4gEHD0i2jKKZxDbjH9oMDnj
Q8FvSx/aTL0JQ8ya0K4xj8X4b02eAbHPmZaGG9Je70TWCrW6ptu0xLJ22eHICAWJ5YXzxyMpvaF9
Qg5iNsmgHDr3rk8sWdVq87Oqjeg+JOzsgOi0M4euBZrAoj5gvn7vDRoSJ4AVHzFfQytT5AaP5QJX
yazi7ylZF4k+ROcZ/YZ7jRrLNmC3Su8TxA5Uy9KOA3Bt2Qr2ijAm1GfK0kz30O/Sm6sn1VIy93D/
6eUGjc2n5AL5RTrg8jliVRX3nc42dnxJBoLw0U2cUBd+iMsvDkkJPps21PmWwDbM2SenRl6GIjI4
o3FHET/BYkC9qPSM1cN3e7AwTzQXMXolUT+RPZbhhY0XlHyFGV9l9p3IloyKPD4dkha+zmoJHlT5
ig1PsJ7rLhPFuFn+aAvgKx8sSjaLAWOfdCZpfZgwZoGLg6m9in9nYQ+wv48oXpZeykzAHWFmddpn
aUyatd0Xm9qjruldGIDdBzdpMKItJa3W5fT9Cy5pJXdrFxh+d13YBwrWlfuQdwGb5hF+Kpr2w6mW
Z0cjArLbgyIEphHyJSI1SGEe1pucHKnOQ8X9npF/PaQeW80p1ZHzTFIqykQeyS5dMfO2eeioSwi6
CDvc8MAiYNYK+AD4tKamHmCWW5bRMVDI6Ig4Ff9NlONCSN4EJjQUJmADsLhXZD/l6S2WdwnShoJx
sOF2iXitGltuR8tqgSmos6mesRkoDu4muOizjdb+V8qLvQ0ktEJB9LCBHknw6Je+QMZ2HB6uNrJm
1wbN/qZwEJgvTXPsSZ6jfuvZ7LURZEEG+XauSuO3hjk0Q21H5brCbLH/fHZ87T+3RgDpGTKgzhs2
xA+dUyPGKgqqccZUyBC3FbM0F52CYCzzFwxdhM13/NafZ11VhCIlnnC8PmFrU4K8QgP9GFIJ9hA7
bxdOC6Fk7wSsMVYIGrBYBqyDgvAj7KiIIOGpI+LFGVFsVkrX+WE9U1YogavlanwoLAczGV7oRQlJ
nv8relbiIdveIQH4iqpOhjLDSlvCmI/XLFy6FCZa+vmtdJJLxRYmtpCn83+9UndWwViovIL0PCBk
a6DLZLHkIu+6/gS/ai99vQCqRqQLlIyFfegrXHsN1wgZGoVoavfbkQfmPvp7DmA/tjwJr+Fblrve
DeIL2x2EtGuQvwpaNy0OEgTyJlidv6qTvnB6twmXaLTNhSu0OJBDnbdA+y7zqejVRf/PVdW5KS6a
Pyl5OdzGcg1UypwPNaKYzn35nc/Wvim0qqx+g5zdtWtywAoh9v/mr1X3mPN3sjCwSJ82CuVzCLHI
hcYSrr2XyRZFN07VQYN2XBSP41wlCPIPIDbkek/AAGRc6IecrNqROHtTNZ2wllSPKrAjA9WquUL2
Gh0daVGWnM5YCptY1BNC+i2C/ChGFTYp9uUbAU0rn6oTCYbyYOY0z+F+Jv+m+zYSCWLpooo3oAaI
6g5HXnUORmssZOqXpCK/ZDvw9fqOIxoSgRpVk2obldsxwRZyjSpijOYuHAqLD1lpKK7oSevy6n77
Dxdvn82jfL2VfUrgXFCZFI9Dsn0Cfys/AttChopYHz4Ba+2FF2lDTZUJqYwzwjYa03DIEGV4r2z8
D+MvzGDM2COm7fiMqa+1WPstqssUYMhx0rKd2i60Au63P3JZ5zEFj8SpFlDZs7K8aTrWhLfmwE8R
DyIGGIcL0VgTPl7vxK1UkhwRNagkpQv89c+dpGXYdMUjdGxdjUCmMk3VAiP+33kjS94hUUzHUNiT
hqTr4p4w/vmJnkayfSEhrP3BECvnMBUh1dTyMGIvPjANXUlPcbGa/PZTFVNW8C4tp1fDVRcO+Ajk
qMAxStg05BUKcuVgXzAQSEbocDdIer2DAngcWgJb30+B5mtK4W6szknCoyYs2Av9+xHcFVERDdXz
vORT6cfKf+5UC5hvOX4LA1aQKHeLxm7wMHPmr8zYFbM71SrJVea+7ovAFDWUPBmrLtmkJmmc/Zfq
LnWum3AsYcE7s30heCFW2kYMHQv84XQNnFOnV8LkF78XMiwwVQGR7EaqRHRxyEiEVyO/ch4AVZNG
uq6ktYPahv1wAw0ZRhOmMvEsA3L9uGZAM+odfntMWtx0XFowVE+jRjPO9vkzsrf3JBgUw2qFPnDw
aalgE6apyYkswt0GkZj3yBmQndzpfP2jp6ixAVHU5McRV6NDwHaNmSkOi6nUsE0EWFJVFj9lyWO/
AuQqPjtkaP1kH3Nhw5JdOCT8vf5TbYreBpAlP3saJi8eUAIrhTx+jsunSatYaaGUkRMaz3tt3AiX
rD0ZaC15FqNbtFobmbpI540xS/cC+aWWYAC47lICzBDjC4sqr/YwyAPKeNAe9oRc6IHUfKeTmWtv
ZUM3qn+xG+AibBA8ULG2D0bBR5doVq4+foCbdw1WtH9aXo9d5JFslNfU6UyTUF/7t3vlCjhBSkt6
bIIvZyBzLXvxJPi5dGnAaDtvZMWro3EKF7qCqx2iyS3TGyDAX3uZbnb2g7nDpSNlKIdaEzssExdo
4ASRzZy/us0tvMFfukUpJzNSDI6+qN5PUkthiiODFTwJp8D/2vx+SUqjUyGaHT4cBCjzW8tMfwy1
hyQ2Fk3rn2QRN2UFWRi8Z/7QiWeDN43NDseax1KZRTgyLZ/s7zlGZLtTxUyXLEuc0syrUtgVBRjY
8wxBm0/Q80K4KTBCud66g6BSZWMtIaJRN4qkQH5U58wHQjhBLC8ZndsBdsR2YoV8jhqtp63Id4XQ
0JJ6/oIf5OWXsrDplXVkHIvDH3icIDLT3W9Cv9p8coXYoLfc7++y309OMZvtLyjQGJzWW+ll/nUs
L5vwtNkEJ3/YbK6jLF9eROjoM8U/uy24n5vcVFudUgK6pN+551A3FR8N8aBHPG/fYf0nNADwgdGs
fekTSVbVlaV301QgcqV6G6uImF1sTkTTM+u34ZLnHQNTR3x/qWEIfLVN2u54b+aI/J45l32kQ3SS
rzk0BZhdHiSMiBC6OOYfhEb40Y/upMB5v9H2N/RrWy2QjwMdGVLp4J4Ww/YwadXunzOIV58tDEoW
tXXkx3tsiBlpa0p2kwjHkSeqVUmC5hIphET9RY9eXXub8iiA1WXUznACdTmSioYr1I2Z65sNLoiT
JmLdLINdflJNTEM9O+Pi7Zg3eTyaQ47g1x5/wsbfuayjm4bhMk3zpu3L881PIYGR/KPRu1BrF/b7
v3MCGl7IYs1Xh+y4bjH3wJ3Hvarx7sFannlB3wfKh2IbdI1oFfakR4abGVZY3YIXj+Xflo5DX1an
y1itrcP8eeCW8ItTQU002wkP+C+SuKW/K8JC68BBDI6JdC9trEGlavXwPTi1/90+ESPVrkfleEei
NwT0SoFsWp/sl/ZCcfVb3crG+2Imfj7jRoDXaHU9zwB0ahZDbmfOpiB2QGsT+xFiek415E9o/LG9
Kt5gaybGbkEkvvgx2qoOtvoia5PaTlGibu3hTTY1JMD+GBH2G1tD0aOQdK5NdxI291Vs0xfA8uIj
39WdWK0Z4tWO0QVd+T3WhvN5x/bk5E8fQ0yhJNxzxPASWwnXQLMcKGIrYz1LV1sKrSmFtkIDEScx
1/ndvydfQIjUUQ6EYOW5aqiwzSKsCj3ub3bSZhqSUr4c4NsYa1IFzRRx5TuYTcH0PmokrjCeloCW
BvmWkF9PYonrAY9uhXR6rFXfDWgixMdE9AVtWWVbLNZ1D9eRMZ4qHb7KmkJ33BvQ3bGPZe2kEcjb
//ksz3FWwdm3XGuYuMsdqtIjgefhWoJTENlYNB3XdqFSVzOKHeUe387TeqbPpzkaTdYXpDZ+otkV
hunKGcbpbRJWycivdCzIzJSRgggTkCaB6MjuMr+0oOS1Uclp+vTK2eWsnxuv8FDy4J/5hP5Y2IO7
zU5nTdYFFBOKSNBy1vmn1VtSJhy45+4pahy6bGe5nxeIo75X2F1oKxRWHQh0g1uF/10u8FJMUm7L
wgtkkIdSgj1kZs/qZUq35HuBHjJGcRqbYfjqgn4Z3evyVTPuK/ycxypypdXp4wjGTALMJG/9/Oxe
ZCzJchEhZVlySQLnuOPK0oCsjm2XG5EamLzlElwbyS/8cmA89RwG0T/+wLnDPQusDR58kX0NOIIM
kj/dEd30sjk1uPfbOgWUqXgKhSZ92mdHMP4YGVQ4Hi7dJGun6xgA80m5bN/7VJdn0Xu9CFm7gu0h
8rxGmUa2b5XCCxbOTjbb/PvQMr5xHO9Hkl/5sUSF1+mWbNfS4njLMNUUh9r8u1k+hqypS3nm4e68
E9cdvoX2ysXh36fO90nmGsD4btA5e/8gKlj3ezF41GZ25QNgOZ3xZX6vBeBCsg6WCluAXhnxWTcR
jBZ82ig7nEIP2N8M4S5bRbBbtySbfhDFP+SwY7ilbQzto6e7axCKY4McB6IkKGxUKoxdl5i+417U
paCZX+og9CndZx7+JA9xUTBk8a/5AMdmsqEybBeqyt5ZtNJDS/1jAcDgoBMuRt0IWnmwxRGawGUB
h6BkPhSNmW/WgGhQ9UqFP3OhKx6vXVNdrTfvGFoSKbbgcmqCDbk8KBOVsAV6RvB1ACZgwACPRUhP
8tmK9+c/R5eqYR6N55cAOn0jG9YOTakoEj3SDNtrke4Lwus+4ufIqVZhOCR0zlkZvafV9HLYLRdD
+m42fpsBnUxlAaUmsnDutaD1ZwbGCEAQTYtbs8den0iasewd7ixOfcZUiVnjGUG0XtsJZj/OpaVh
s62I+rt1Ev5uDpAYqVnc8s3h2/Z4uH0e9J2oiJo22ctQKf9wQN35SsQHJadLpQhfyU298kxiTxdh
ul9QjOEMAGLcbTkhxQM4VwnIVBgqeByeZDDsqDm2QSEf0bMNqhw6OyZK40Pft/aqQBq4Yd5KLNUw
a4IxOpY4xM+QQjOdYRCGBZ2oqTKKCL/lHYpHE0A=
`pragma protect end_protected
