��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�>	��h��H~,
�z�*�M(�b	������LV�laD=tp8F�)	�ŀ)v�ޑ"^��F��L�> Ó�����M4G�h�.Yv~��f�+�E�9�?���;�Ω0�4��H�;uS%."q��Zd�/�]�+G|��Ԇբ�n�<!�?�a,��5_��=�n�����~t��^}��ٸ�/��eLУvi�i���m�ޮ%G����i�}	�71\&��cq����+�zE��<�`\�L^�e�|�ی�k��=OV�B�v�@�1�^'盾�R��9��'E�򛚤�p�E^΂�Ok��������aG|#�	[m���}�����R��=��ئ4�r-����[�}�x� �|�LW!�c\j��:���ȳ�oi����_v����jqQ�#�d^��Fџ��<0�
)ߪw�B��ֺo\�s)��M�[��	�h_*9o��E_���]��F~�#?ٌp�&�5d1�)G+��� �n���?z!H��x8��U2�#��#T�I�%j=�մ� �Q��9n��C�)��Y���h2�'����lw��9\7�� �9�`�ꌗe��c^E���2;�%�R��� �w�Pk����9���sr~P����u|&��S�-�}	%N��v��	T)%O̘z#i!_ ���*�w�3�Ļ4�L�~�Ǌ���R�o��%!��V��R�����	+ښu�u��a� b� �$ɓ���������G��*�N�
?A}��02��߫w�<s�O������!&v��šc�lA��&���h�"@$��H��r�l�f)��b8�ۘ7c ���|�(<�1��Yh������*�㋽.L��E0pa'E���d�0E�J���G�?�X��$�fxo�#5�P}����,����w��g�VN�V
�#HȎ��U���̏��;Y��c4�p�C��Y9�\v	�5�MX��Ǌ��%�1��9x��X���Zk���j2 �5)e�-oO�P�]�ѐ��n���F�T����
)�@�s��t�P�܆�,\F�Ehi1�������"W�_e�y�ͦ�>>~�/��};�Ӈ�1�GҢ�m�����
 \ n���&��z��e��� ԺU��欀�Iv��ow;�V��\�}I��3,j�$��	�J> NF����'�	.�0����е���F�Q��]���c��4~�yڗ�n��⇩��Jd����v�ѯ�3��(U��h$:�����[���L�&����8�}��,E�<x2
ogqҶҧ��g�ɸ&c��� ���~�+�W�u�(����fK[���s�ۉ"�Yޅ�f"�l3��0) �C6��srV���0��K�E7�߱��lz*�@��:�m�zpX��hFmx�l鶆F���-yVkײ����Q��[�ZEf�)i�OdT�A��c��
���g%�j����7K���1|)�[�E�$��	269�����U�!��m���
��[gڬ�B49��/=.	��+�)t$7����t�6��$ ʵU��伄��w�.G��I����^<q'�A���@+h�f�V�0���E��:�GaL���m��MО�Ͼ7=��rO�s�A&3���e,j���[��aR5�ô��>�Oڦۍ!)t�'W�C��Lu��w�@���PS{+��������Ea'ߒ	�]
��8U3(�?��N�4D��sOڸ�D٘Q����slI�pXҷO�n��-�a��̡���8`�#,C:��3���Jt/��m����$ڽ�`�q�Y�HÂKl�
���2C�Wz��u�=9k\�b�u�s?�(�Q����>��-F�e�O���Qn/zrD�cؑ@��8� �a��4ۇ?[�l���kL�Y\�+���&��!~NM���(�c��m`��H��+�/{�ѝ����hBJ�����Nf=�.�pP�jc_�����Lɚ6��q��|Q����6�]��n��H+�]iʓ/HtW�?^��_��	`����]��RS����t�7s��<>��J�&���c#p�{ɗY3�BT�9�.�Aw�y�<�Ʋ��k��e-����<m�'�m'1ZV��_�)<�	�*!*�L�c�sZJ)=��^n�0��	3��K�T�~�1|?�դ�?�E�H�����HO��9��(܉��/C�JN$�{n�w%y��0Z`ѸȠP-#���}}�__M��ɣ�E�����MT��� Uy����'TY���}�PN�u�������N��]b���ݶ2��L�LyO�w
��G����j"�����6=�i��h�n]��*?.p�?'�#�L�O��K�����c����L�"Z���_9��<T�h�u�8+����)Y��<��C�z���L��P�)|Z�|%���9^iK�����q�5K�������&���m��K, �_f�젗�0���-:_w-v�byZY�5_�E���m) ŷô?u[ٌ	���ڼI�-�IX���ϫj;���u�ưC^��4��YS�����VPcxX�6$4������Tz_x8�B�f�m�==�V��D�E�|SQ�6�oN�m�YԢ���Zd�����7 �yd-a�J�iPZ��6N�Q��YP2Ǹ}[Cy��5�.F��L�}�����ݘg��M�+ U03:�(�o����(��w��z��WǨl�*��t2�,�B�`K��,��8�e�o�3r�$��=���#e�$Z�WMK=�L��l,Ub����61��	�Aϊ��s�<B+�tD*N������B\7&�o��&q���6�Rٽ�c��[��<�q>Z�/�,+�}p��s:o1SĢ{�ω@1��;�<`
j�Gm6��B�s��2g^+��I�����*-j�� ��̅ �C&2��nR�u渿@��ў���� o�r��#Q���*��+�,�~Ѓh`%J���!�,�'��ڵZ��B+�/��d
ab�"S�-W0�<@�o�������pލ�2��:�?z w�8 g F�L��K���G�,	�"��\>��^gC�
�=t0�޽�ܡTT�^85����t�M�s/fئꞋ�8O����#A�)L�?�j�m��|��oH5O5 ~�i[b��j"m���xD����Gʨ�����]#���Oٯ���˄�$�w�U_.&R���	gc��̉��m)g�8��SaH)�5)���v̕)���.��_ܬ
u�o��y�=메�������>{!8tЁ|JΙ�:n��ҙ�2!'[�����^S��:��w'�����\���X�@~asXo|�kGA%���k;���s�e�Ճ�MZ&H���BpM��
�����:v�}>��`=+\�O.yw�]��K]��1IA�]^Y+V��U4EvB�,;\Res��W��0}��5��z�-��u�I�"Ee�S�������;G���a���b��z�ć���0
lȶ��y��T�T�$����S�|F�q�@�E�R�a�_Ԃ}�İ� n��z�5����'���ų��!���^�Z�N2y��ZEiP��q °��]�ڍur��g���`ci��!~uw��8b�8����D���A�sj|��D(�cs}.ꂶ����
-�n�Q?,���s{sY�|J���s#�g#,��I6od�5�4�89�g~M�*N|���vm���<�⌔?q�->�X�5�ٲ$�NN����F�`�������FTj(?��ؕW9/��A���o 
PnS��2j��@DSA �
�擈���U\4!�Rn��op��y�t'�'=�lu����ӑ{���r?f"����7`�L1�rTy9l��?m�6*�i��R��d����Qr�IK�e���r��Ø�j��?�?<=��<�O�*k|����.v=����8Yq����S�J{7Q�1/�;�7�ڧI�#%�AUu�I��%I��>W?�O�o�`��'ń�U�Yy�	��rwZO�.>�~����}��b#\����o��=y���؊^� </oN<a�F�X�^�L11~��|zz(��[٠���ȁ}{��\�/_�"��O�pW8[�S��@��qH�O}�B�L�l%{�V��l��Y�:��ϣMz���#Ơ�]���p��������[���$��w�ڼd)h*�w<Ů��$�3\/�?���C��"Idc�}�w�}�&#�4��s��� 2�޳%ҿ��Ueo.��i]iC��/0����m]xʕ�{�x�+n)˃��.��2�cs����m�]?�4�.<l~󾰍o,��dʖ�I�ݞ
�9Ӆ��${��|
�{.��q���\!��T<���7�D���]N�+�j}�_��/e�:%�we��^�_-=i�Rl�&X�H����¹S�5����q�N?U�Q��}6��!.~a@��#]��x����\*Y�%�-	�МQW1.�l ��R5k��
�0ޚ�>��r�o-~O�i9�� i�$����W������h����g\(}Q��&�l�9N�WF���ֵ����.��?u7�n�CS,�|���0�wC�w/=����y-�*�N�
*���)wc֚����7����f��+h,5Ɔ�����D�0�j�Q�#���ؼpG�Q�����%Ci�[UVle�г�>��Fj̳��;9=<��<��A;��9����rP�R��5���M���������b͵�(�1���
�TZ���(y�߳� ���N5�;���^�GT�v���GG��q���c�A�E�WS�Oe������7bO�����ߘ!�ORqe�w3������������n5�sK	�?;%WF|o��|=�%�w��tp�M|�:%��H���%Al�{,y�zYj(y��k�է��4b>k$�YLC@���ቱ�7A�'��e���i��8g�ø�梅������b��	N����DE�S�����V�`<���p����tY�yhm#A~-ߎ���1�"Qr���`/5n%��Ǵ��/��Ћ�OHeY�s�O�
(�Hh. ����8�Mҍ��l.����0Q�����p"#�v�:D��<�y0�t�,�$c�յ����~�G��{�J��I� "����g�Y��cB�q�����nƝ��8��e�h�'.� �/Ws����u��I�(�q��wM7	��ta:�<xT(�.>�	����gb�pF��+9�&��OHq�c-�|���x����	<�Bl�r%c5&>:ݔ^6��@�$�����L�|q
�W1�~C�Wq�+�0X!R4�0�n�O�6�A3��~Y�a�B4Q�A�u�箑�I|��^7b[S��<dG���tϽV�K� �4{[��~��b���p���	��ي�n�*�ɫHf��.��:�KI��~v�Nr��F�9�CB����;�U�#�M� ?�ӹѧ��\�j��4M�����3u%�[�y���8��Wq�\V�C-!��ui�L���O�c�X���[��������V-�:SY]&.�č<�#�n�enDR�f��x �R�F;Z?HcXB
�D=���!�l�g�C[��>4�Ft�%��f]��A	8ka0�=��8-�2�9@1�r�?����V��y�SG;|��@@襉�0?�V����FwK*���Ӵ\(�@��ܖ ���U?m�Td�t��ϴ/�Qt�Ua�E<��dc�E9�,h��ty���B������{���<}leBխ��0o���E:w���U���@�j�W�Ve0�q�W��vd���]�̫��''��[6����꽯��J�}H+�YĤziTe.��-�8z�#)����H�� !�үl�Fh;ɾ��"���'&�y���E�= �o]N�lVm�M~��ݷ����@r<qTG��r�:hʞ��I4F�,�TeB�Rc�����qMX�YORy��E@H��EU�cLE��� �A�
:��eT��x� �b:g2Y��;&�Z���J��[@�9����r��"E(e��]&��6�N6�dSx��P�C�J^w�F�t<ϫ�-�(JJ�}W�ܤl� D}��=>�AS��?t�ջE��\�&�ɨ���`8|��6@�Kd<��ę��A�4nې����'�+���$@w�q��#S��݁9�0��X^�ܴ�����g�8��2'9��Vu����BIۣk����%%�=��1��;�¡qV��^����⡾��&9��S��]M����k�����T���
��#D������φo��`�l��Ȧ�0Kx�+�ՉOSQif�eNӶ�խ�@-�q����b)�����*/���.����H��Q�1N�'W��E�Z_a����� m_�-�U���DH��Aȱ��b��J�v��0ʹҢ0��U�댸�M���f������3��N���	�i���/���n�[�(�t�Dbuu��X=PZ7�D�ѝxr�?��L����E��_r�L�O��&��*DX��U����Q����x���U�9����X�(?=�,Z��r�d�X*(�)s���q�ɂ����Dғ��J
�'=QLh15�$�V�HO���L�[̰��qk��X[����e㝦��)K�+�m|�[,1����`�\0��H�L�簺��m�����I�c�:�{�auF��!O��ơ`xHh��Q��^j��'L�&����|���S�-Yպ�C�'�fb��a>?K�c�H�f��ě�r2c��# ��ܝ�kx���E�z)��.ޠao�r[���̵UD E���;�6������*��ϯZ�T�Qm����ėuF/ۮK��@�v�4��9e(g��i��$��d8��]������e�^2$����aX�r�U	�-")4�����qE}fx_4�+�A�����`�]�p�#z2������vv�X�Г>�`0�o⅀�-�w8��y Kb$מ����0NT� �!��E�!�9�U���&JT9e/���/-\�_����I��j%��Oh��TZ���|u��]*��NB�V1G۫���~G {���E�{��E�n�L��@���{ya��ٽ�_�e�.��jt>���+J샯�5*[�j�X~�vzx8!�e���+	��@ȟݡ�	[�25p���U���	��8���ws��c{�c�I�л��4la&lr������Kh�?$qv�S_AU'g@�v�)m�;!.�6�|_aX�o����zSM�~�d��Wf����^��|p�]-��NUo��
$���rbW^0�ַt$��뛕c�?ʾzg�(l�}��٨��1Ne��Ymvq���z�X�Y��y�d}۹��#�~_�3�P3B�]���p�*g�\�e�גRĠyוV$��m��`�K,��迷��W�Pw�W1
�� e��]��C3cН�������k�+��K�:z�U��.��!� ��v��Ψ�Su�kW2U5��,����y��1��*�bn9�:r�?>�Y����P��[�%���6��G�5T+4{8<�u�9/q(l��\J؉���$��u�詐��b�Zn����@��E�N�F���6���=�!��5*����htB��� ->���_e~�i㚻� ���]��Id�?�-i�P�qӮ���=�=��1��$hmw��Y�K]��n��"x6�!�ȟk���i@?۪g�3�)��<���D�.�҆���@#\�d��8����}���Q���k�E�=�I�4��2�z���
�}<I��7L:��6�*F<}O���p��ϭO�2��թ�c�̇ad�^�r&�d&5J������&������9�p]�t�B-�S8�4�"�"������C��]��OE�MPPk<뢤�4}=^���E�S�t�8������N>�wd!f�S���q}����r���;P9/�9��ĦSlo��ⵀ5;�y�m�x#� ���jެ��א.Uq��w���.����v�L�)%/�{�F�Kb4�M�}Cc�!��sU;��4���H���&�,��CujH5�:�8�.D t&�^��Q�'żkJ��4�z��{D�L��+}S͉5hW�����Cs�M^ �����<���C�h����b�jq�J�J��,�}K�8�,�T�[�'�ƃ�IN�.�c���6\ߛB��ғK�͘9�x�'s�~nZ{~��p�U6i��5���[k�ؤW[xE�@��C��&Mi�xV���4�ҼO[���i�|��983�F���|{U޸� =N���1�e^��
���	�"1�����~�ٞ��o�@�n�)Cа���z�~7��9Y	3$��k$k�����Ϲ�z�7~ߔ�$m6�11�"��̋�1������u�%	Q��MZ�Q8���(�i��:�L��V�E������4o�/��K�aG;�8A7��E:d4g�oE��$&jqY���e�P�-���h,Vk�}�V��ER�e�f�;dW[�Q�)�B*+r=�̵l� �?Dud��nĀ�ӣ�+4(�O��J����Pn;��oI��A��;f�e�r�������2�0D`}a�KJ���� �|z�DZ�]g��5�������S�A�in��0��9B� ei-x�c�Wx�e*�#�+V���Ko����b	�Q/���l'���tZ�u�3+@��a\�c傿�E���A�?�]��z�96j����"N��e��X�N���>���<�@P�Ѣ��QX�I~��z��K���=�5�E~�m�'j6gP�<�$��� Σ��߮�`;���%Cxu�՘��.	 ��ՙ���V�i]�t7�Tᙘ9�3R��Tђ��_���%�%X#��0+����[��^��Q��w_���`�q���I-��d�	��\Hg,��X���;�Yw��t�Ѡǔ����5W�ޕף�c��g{e�p�n��lĿ73�l�eDi�m�S>We���6x����hE���x��?�g��f���h#��ڲ j˓Nx r ]���t��z57�5�: �ٮO��ˌz��C���ˀ�K����jƘ���&���S�q�\�A,)$gި��9w�@�`�w�xz�μ�ґ3��!�(��#���W[��vW9�S*���W�.��A���{1m.Km�Pk_l�@���/��|	��:2�9z'i��Y�)2��&s�fhl����cݩ��{��ܲ�V�Ň�^�?�Q�?23�> ��j3X�6\w��V���M����?�,��2�"rB uTo�P�*�Bk�KoRa7��D2�;�ʃsqWХ�zԱܜw�Jp�/NV�	-8S�Թ��;��t�Z�[�$ ���^�v��̣/�r/8+������T�w��DU��R�(
]A�}kn7��x�&(��:YZ��y�ްԒ[�~�*_�e�_���.�2b�0����G�7���W&�k�Z+�<�?�Hw��E�E��6;�mx��M_�|�n����Dg�o�<��"޸bT)wu�b;�PyE:]�5Q��U$�eϦ���bк�J����3�?��#HdX��0jՠ�s)�ŒTc8�ڤB�,j��Jv�[�6M(Ə����"D���e.1⢌�Ї����o?�@[F?Oow��ϗ�/����<��
�m��o0�� f:��9
f"9l&*憫���H2�W	 �o��DC �<oX�5*���U������A"��}1:��ys�!�ʅT��j�k�lfj����2��o@{�[k�V��-�#".�b�1�]���w�>bգ�xޚp�asH܊��\�.[��Z��{$�&�D�֢��4s��m:����\�3�r����w�Q�P/�ؘ�66�Ѱߗ�*����À��_ɩd?�����H��]�Rd}o�U�m��ZP3ȱ����H�C�!�:���	`C�¶7�q���W!����K!jwl|_�?�$���?~NI���T���K��;�oK�������Ѡ�Po\q2Z9��Nk��0��]ECS͊�Bz}/6��r�d�v�{F�j_'0,��%�r�Su3��j�C�~/�4	1�1��Lu�<Bf�Trp�fW�����R�­��4"݃*�rj�t=w�wU�4C[��*r�!1_e�� �yi�!�2Cy�^!=�<�Pj�62پ�/u���N��5&��9�hǵ �/r�J�n�on�vQϳ�w�<%��u!Fi��<��J��
��q395�1QI���i��E=�>�
�r�½�����-�-�Q�w�ri�ؚ��I��xND�5�����
kX��Z�b��p���q鞠.2��H��o�U�z��}ѧM��T%�����1�'cl�J�s2��t\Io��j�����r��Y���F�/�Lc�Q�⺁�{k��rOxInsԽ�.��{<�,1G`R�����y��w֕S�䥹[V�X�󚲥���O��׵ӆ��~�����.
Yϼ�~|��WC���-�l�K�h⢋�rw��c�T��|JtG�~�k���u-/���$�f̆���X�*W��7@�bU���8j���Km]4�t�D������Zd� H�3�,"k���u6�N6�O�W}I)�b��o���L��#��G��|+�\��{���g�CDּe���i�c>YH'D�)(��P�͏Ȭ��!zYojǹ�P�N�����u;�avix(
"�������K�,)h0�@f���E�<����A1CS�$y��(PH��? (LZQ��%���ͳ��$}MhxUo���Pޫǆ箎�;����f.z�
a�~��_���v���Rp�f-�R��\�ls�*�\�� Q-��ݟ5���YpkY/*�I#\�l���AկI��GU�`f��fUj%�n���$����4^+�Vc�y$��(�؇���/�/v�7>�s�����V�5����:���~���{Ô��2|���W6�r)���c�~�v�� ��/�3`-y�@�}_ݿ�C7�Z����4�5��{�M�#�X��1uq�U&%�cbH"����p�&@�a1pE/��F9)I�TԹ��>�|�[�&�̷m���u{���8�g�C=�\�?:���E��ws���So�ŖH�0���q#��ϗ�Ԉ?M4~%"^�@*P�
��,�@�f�w^��l����v�=o`�EJ��l9!�.�Q��]������ϱ��U�����m0R��>�+lt)���z��QTP��2���8��'m�#�\��G�g��0<����f�.�?;�x�����{�����m���gB���W�N�O����2��ifvR�:W��*}��5�d`@O�Ž=fcm�j�J�`q���'�r�ǰ�Lw�-LN�i�m�
�k����ƐW� &�\:f��ۮ�Ņ�djS2I㸘�+$�	�;�a�&�j��7����X���J%2�:��%���R�� SV&�.��+2j��Ҫ-�IA�`��~��w��;z�!,[>|�h�[�I��,�z�
A H=�_֞1㠚������ȁ!�FT^2K�)w79+vrD�ʝ�A�8q��q�ʀd(>�41e�Z&i)n��a�J%s�3'�\�	��,~o�ܝ>7J�~o��k�ڢO��-��ίne�-��2j��u>��B#�l���p
ޅ%e�xg�mm�@��Mj��p*�[i�,��;�v���q��ؓ�h��e�fDŵi�ތ�S�r�d�v��Z��Q̧�"�n|��BeAS^ٱ���q
E�oM�_�#Pf�\xp8�����w�nD�0*�J|Y�	ieK�����֙�1yUt�`a�0��̹͝��$[�6.r�b-伮������������V����ӄ_~�~�0{4�nw{�>���,B|(~��,_r�
sˮ�\�*BS�ݪ�h�Z��Ӟ�����+{2��,'�٫ڿ��yˇ�t� �S��!�� e��6V1ʿ2 A�����6���w���⌛G9N�����yjKzav��+X%護�)������#�`E�"�^|��#��e�G�h�K�,$���
b�����5>;�V���f��\�jc+�����Xjф������EZTr��,�`�����x�Q�18��L�[\Ƽ�L~�u�(!zt#��=��RȆ�K��~e�!k�Jy���3�=�Y�i1�
:�ͭ+u��m-!'�N����c��m���W�=n����o>O��ݗ�z�D=�����m	G�����+p�������z�W�<�AwK*��q3��gga>2���|M��<��$f@!y9��z+w�N1��!�m���x�(��K��]�.��T�����c���s�'�c
�w�P�C�|��ؙz�1{�<��WS2�v���)�|�=��X�DW79�e?Q�͎�!)��s������֠4�$j��D��՝�J�T:�h1�"���p����p�Y0�4���2�:wA������ӛ��'�'�#�:�����Uy%��E��
�ţS�U�sr� 8�G[�'��8��Z�@��
hJV��A�mp����0�b��S���i�o��F��A&&/nN����􎌌�¢`�;��53���1n�꠰��3�r���6>;����>�T�r�Ӿ��D���m���Ɂ&1�c�T��:3;��#G����Z+�i���^!��2����h�_y0R��������"A"*����XbhH��g��8���*���ֺ����'50*����xd����f�b�~A����Ծ`��P�Yͽ�]��������>���l�bk�lh��Q�M/��+\ߠy��ҽ�c�hb���3+�h���'p�#�0����()�$��)�b��Q���y@A�bS[;���Du=��D�IQX��L� �ʡޒ5%2���/Q�����gZ�����)M3hjǗ���U�j	��q��ݹ���
@�4Ƌ�O���^p�9:��fS��fຆ��Ԭ���E:�;<���ǝ��W���.ݕ�s��Hߢgc|�X��!�{���W7�!��3v�3Te��;W,:��ٵ�xn����hO�t��,b� O,ú�B���.V���_��)ѹ���iƨa������<���^��~C��l��!p�[zɃ��Ea�bϴ+u{��i����ג��{O��`�cn�^��G���T�\9g��y�\N�����Y�3���$w^��\�t�N���MU���6�x=ܘ��jg��X?��TKCw��h[�0�!�׫DL�#���<�{��g���D�g�Ѻ�6�O��.5V dgu�$�p3]�De㘐�t� �	��|�Qb#��h�f��Fw*�y�V�Q�K,)���}X����cXl���n��F$�E|����[bh������p<:~�X0��j�9]ez�0���7�nxU�f�#�ۙ(<���@V��tÆ�3����U���AY��{�*�����UI�ϵ��b�>���
�bͷ~��ʴ8�! ��6̱�FJ�ǟhEM���\����/��\O73�2;��#h]��?)Ig��w����!��0��Wh=��O�pn��JeD5;a~V���j�G�W�a��soW���g^U���{&#1"o8�=w�Zd""h����w���zI��������f�L������Nf[�g��^ SGU�o�$Dx��rB��_���}�����
]t[1�ñib7�K�-�T�q���u��<_QJ��O��PGj��>d����{"�D�S��d��YK �������)ej���:S7�>�I�g��m���xT��N��(bb����D4A�(zd��N��:�0�p�۹������uh<�d%3�l����W)M"������cH`�~���v��{b"�[��< �Xp�D�g��1p-mk����O���$�=5��0mEgJ�bϑr��T�:�]{hR/Ӝ1��9 �͐�nx��+��G�hy���M7g�6�b�Q�KX�4!!�U��e�xs�N�"����R��	Sծ�GM�ydH��u,�QZr� �~X�P��6�l=�d)DʬQOWa�o��� ե)�[�m�h�϶J�&�Eu�%�ۼg4�sҷ,-���,Q�W�u�gI]tJH{��x�B�vF��ʨX-r�̜.�� ��F�z��p��I'Y*�v8�}�P�h�X0�}��D��d��vi���hi A�"�i��=�N�Zz���_���B�^L������q�.3�i� ���������~Ֆ�ǖ �ŒաwW�`��uw�^M�p]����9�f��Wz��C���2�j)�uRɉ�b����Kx�R={M�����6љ�����1k�u�+p��m�[j�]�!��a�l���F��,.�s�L��JƏ����if�NPyU �S�S�T�f�Pn�˱�Z�w�S�,�e���0H&���s��I��9��e�Q�h/TɃB�*�	�5���N�� 95<jaֆ#�w�Û�I�᥅�B%ɁsXuI��O��X�Aj݋+���=xW$oG�y���T7գZ�?��6(�LM��f?I+Cl�ju!�O�o�.F����6�Bmo$��!�ԁ����) ���Vk�O��1u��:~�EOK>�:b'|9� �D�u�],¥�C|b��ov�h��#�!�g�;*ԡ��Q����r�1�<&�|k��ph���oȇ>�;���U�}�� �VЯf�c���̿��]�~����Z)��ɏ��\E�G��{Y��!~�2��)�|���0�H��)Ƴ�HI����|M�A�7ݘ�XP�lB�W��<��nCCtQ�j����c6����;[hO���h��!����`Nv&�j�!^ahŇ�[�XFkd���Lz������Ugg��}}`Mزr���`���ꏹ����������
G���5L�����.$Q���i� ���3ǙF�R9 "��6!.��Y,Ȕ� �R�6�Y5�<hP-�p~HEI\>��X���f������FK���Cu�".�q6�̄O��A�{M�]�LNc�9��P�����
�أ�4�B|�TD��W1��"�
t��_�f����ţu�������(gn��������� ��ҕ�}�"P�%��u<�F�̠ԸK�h)\`в�ēH�B2�1W����i�-�?R���s=��KHM��Z��f\���7��jjCP�w���n��M�a�#�u.�f� :�kz7%�G6����H2��l�3���}�<�p.1�E����/[>�>�-֛?v-������z�W]'r�(B3)�.1{��Ow�(�@���h�ۑ���A���[��� ������o���EU��P��r]�g�=��i�Ps�GǃZ�������ّd��rC�"�)ߜ��q�V�DgC��F�IGqc�Z�_���|˸��kt"A堾�f�%s~�s�fQ�BK�j>�%F��ޡc�&EDJ�񓚁$M���~>��kw��_�moܿ[N)+��w>:�[�a)=m�W�&�M�X{H����R<WG�?�Y;WfD-�b~-ܰk��O�k��u�(�|޿�l���a�&�&z���X��2���s�>�"��	���$!)�Xz�'��*%MG�SK�`(�ל�yv��Y�m�k�U����YX'fQ����JTqWCxa7�*٦!K^��R"/Ki�/�,	������r��*���N��̸�7{y�ᓧY���[����p��kh�1�R��L��ж�q���6v�����N��u�џ$D�P:�0K��r����r�}Bh)��4���M?-k���O����-r�P�2&8���A!w�;�#�}�3t��Ћ�,%`I*ʷ�!"�ضel�^�^7'M�`�
L�Ql^kf��������rP��(e$0�����*�<�Jlu1�l�b�.:��@x5!_2?��A�!#}J(�paj���Q��ULL	)A��Q#�Ж W�������{��i;B(���MH���y��6\e��G�;�C2̣z&u��|���K�h^2��NW	w8��Fx9Jj�it@�s�a�A5�����z�mz6?������2m"+@{8���Kx)�;���`W8�`�Zf�A�L�\�"1w2�5���K�j�:�t�o|�lx�=d��?�\�|*���l����s{� W��mn�D��%�O��4�HŞ8���&��v@#g��!�;N���cE����9Iz�ؼ��Z�)�� ڔ/��bJt����֚/5ss¹� G�A$;g_�N�8���#��Oh��{ �wCk��x��m匸w6D�+4%�yyM�<�S��WHH�C�2�߱=�k~��rt�i�ûQO�D�Cf��,6���-vj�[�B���E�D81?XЮItgon�A���kc�U�F���˫3���'���{/@ �\�G*�檥O�M��r^/�C�l c[ź�..R�� �,�Mv���i �|��s�2�'���|�׶W|��[�Bb�/� ͽi���	Tq]V��U��[ߌ�z�(�t�� C	�F7���R�K6@��=R�١ѹW���7��k�%���iU��N�8
`��r�VNܷ(�����K�ai!"K�SHQ�]�pV	W��,T����+�o�	y�H�\�^��'�a6j͗e5S|_���uL_�-�MT,����L���_]����ȏ��\�f�p2s�:��x
���:��V��:"}c�����z�����@���x���A�~�:�C����J$J�����G�X���3�ܐ�ݫpMֳw�ni8��R���M�- �<�r�s�0U�Y��V�%�f��ND�齿z���**��c�_ϒ����Y?W���1L=�s�gg�4K���>�
F/��ͺZ*�{���g{��ھcAk�qhYx�d��tkt^�I��I@���������}���N���G�ih�_��w���~�a'ա��|�_� �]cl�� �\�E��orܩ�H~�Uޖ�M��^��x#�y�E�*�
�FZ�Ӈ��q82'"9gj��J�h]�gۭdo�t�w,3��uj�U2e�d ��ؿ�7������O�n|�1�TD�
<]d�9�����\z?�1\�9s��~i�dW�FB�(�90)���l�k�/x�Q�F�GV��:���T���N�˶@�7�F9��ʣLP�jo17�S���&��v�쉓�7҆2O!�u���&��N�	�>��5	�L���{6L��#Gy��KS��3��E�����HS��`�a5�(,��I
E Kn�'f5*�;�����wc�B���Z������B|%���A��`a�i���P��'�zk�=�Eq?��K�Ʌ�/O�Q�n��I���sԁ�nn�Zi- ���(j��^1q�����g�-�����$w��Ӗ�_4����@^]�߃<����L��G9����a>]#���oD�%�ݠ��:��%�;��D��`�A�`YO��m�=m�`,u�~dŭ���.E�47��cV������b����f���
��Ҋ�<x;i�H�2r���R��(�@��$[�>�AN�C
a=AOs�聳:9�YE��x`c�A�+=��\7�>�5�� ��%�x��n�\��������)�%�?�!%R�W/�Y�n0��
q�����M<;*{K"u8y�>~5�|�����4`�l����Z$��5��}���-��<���ɂ��*��N⋌f#�gi߼^Z�v��G��I�F���Q���z�=5�)�����t�I�A�ǩudz���c��b?L��҂"�JD����>���W�^I}������oWK�1��#G)�K�࢝�S�Ho>J�� u`߻d^�njK=��SA�,��\�q�`T@��ʟ���Y�gK�P�S.x2�v�/�<�w�V�͸����b�*w�Aȹ-Z��+���R��w�P�F��u5U�f�2�M��}�N�ad�w��N5�k3.7 \kB�_�Pl��y#���hq��p��w%�Y`4�u4��$F��bĉ���~�lX���|���
�<q1���|�@�j����f��}���6Hv(�.�^*M7�
�u���*�T]�`]�(�_����C�� ����_�Bf}�څ��9���H����NڱR�/��c~�أ)�I_���`_���ar�{A�:� =J�{̃Q�*�`�E-���l�j��ݷMͦ�>��U-�I�$1Q��ywv�޵��F�6Z�{��q���tO�����oM��G��$�T�6��uwv}u;���8�`�=RF�������xl������:��g�l�s��!�r���=���ԑZspݯ��0�@<���?��b���⇩0������:��\����T����x'P�qc��z��]�1Ԣm�8$�glcCMMJ@��;����#,מD�48|�њ��%��[�%��%@��Z=xn�<�w�|�̬��9ؠ-�Z�쇕�_@��u����F���!��Ɛ�$D(Qd�%���
$��lW�ȳj]F�C��Ȏ�E��D�Rx�S�IR�������{��硝1\�l��n�s�mzIA�~WǬ���é6�R"d��"��f���~��4VC�X&���=��B2.����%����$���Z��
�s�.����D����`�W*C�#�l8汳���� ����3s1�|/��`[����0U��ׄާD}�L�2�L�p����y�Ty�:��xh�����螩[vS��	da��*��@z�������d��}đh��Ur�.�A�m����ì6��=���a@=xN��z��U("�[���7Y��"�KJ7Ҵm`��oT������<L�^V��B����(Fv���_��p�z�5�ٓk�I�%��������;��[�b$�j�tl=j�~N#�٦<����ǽ�8���;���%�����/DV��+u{C�X6i������d�銡�\�OHY��2�˽�E٘��?��ż
����J|:���ޓ��\�SmgL$߹P���t���q����5adE!@C����;CSMr˘��3��
�kSE����=س�X<!8����Ȱ�����sE;��7�Rc��4uF���>�#rNeպ�u���W�i���h�A��d���[#g�lh��󯬜�X����J[�����Ɯ1�~�_ ��[�RG"��C����-��b�M'-!,g!Xu!B���ՅuBq��=V��Ӗ��F���Y�(M�4��g��P�Vdq*��
�90��^e�c+$���F$��c�,�L�I�|G��>-�P�w���wJrp�=���OU�H��;�!^$���Lz/�U\���"w��<[�����4��"�Mo�z:�������kE!�~�;Fߢ,��ٝ>�@w)�%9�4
�&ƭL�m��~x���� �(�;�rl$W���f��_��XN��5�n�S"�.���><Y�t.�l{Jˍ����,.�ߢR쬶�$+;��O� �+�t�@������t����;�+�\Y7�}۝x�A>��$��O���X��`�Ŀ��z��
KN���`v2�$q���$a*T�U��p�?���.X@Y��P�e�P�]23H�|����v��m�����;�	���|���%s2�t�q�m.��F��8�J�ÒT����"��ŭ'q�g��gL(i5䤊�'CB�2�A�t�S�e�ɲ&��K'�$�">.���Ē=\iT���%��������s�.��{q���!��e�rY~�֩�y�*2�s����G�]��@�MΥs@c�#��jazI���]�T?����2H�J��:oa��z���{�u��i�٘��c[�B������C@���	ɠ�l�57��M��ފ(��p{ ok?��&K=DZ�⺌qBt�a؏����V��7�T����k�t�wE��\B�C�ŕI���}2������B�M)�\�VƁ�Tn�^Jr`��I�C�t��l�w����t����Rn[5n`O ���ƪ<��y�_����w��t��5��q�^�٦�0�,Ŷ�2Q�YW�V*�����Aì ��1�rؒ�pBq��=k��=�*fk�I�Hj����k��c�s�6�V�a�1�wsR�V�3����t�?o!s���_YB�~ʛ��2-�� ,���� ~�;7=l���4k����v�0O.�g�.�,�
L���w|_A�퀕j,d�?.� �o���U:���ޞ���t�����R�V$)�-��k��HE�k��Ƒ��w�j5q��B�[�OYd��t���-�>_Vh��4{Q���Ւ���}�_]�b[�+/�~�u�>���*�r�G�͎nS@<$�1�E�B���O�Q7�WаǷ�|�]EUv/Xg0���6�&?�jƹ�#3�=Rc��Xe���*CY��S%1�Eqֻ��Țl�jG$��;$�ٖ]m��>��0�g|��㗵W�"�����g1�����bD�F�7���c���G��v3��[G��6�'b��7��݌�q�z Q��F�T��r!⃏d�pW���<ųj�3dhI�.�b;��q��r�UU-yv�XΈ9�T��8�7%2�Q�,���'\Cv �{$��G�j�9}�_}�������(ZI��
%O���B�P��A	��א�!�V�D�x�*��g&n>�=����̐Q�g{�&O��I���?"�IoZy1�"T��A�7N˞��R8��s=���,Aݜ]� ��䓟��?���d�M��/�e�E
�{ҩw�>�F�
��F[0��j7jtW�圵�v�@��!{z�;��Z�Z�oG�N����ȭ����C?��r����T�q�IxB���>˻�Wy��e�2gA�F�F�Q�K �9��l�������(:�D5b&��\i��p{D*|��nx���S��[�'�l���1DN=*='[�8�)aTd_�ބ	6�g��2���I��`�2q�����Ȍ�v6��t,v�K�(mU(�%�zD��ftL]1�#��˖'姹��s�07Y䭑p\ؼ0:_q��g�]5�_�*��D㰖�;���m��g&���sp��˅WT��m\�
��
-���ٝR}�L�;~��s;�ɚ3O���P�{>���+DȆj�J��ћK>�ׯ&^�]�ؐM�\�A)�6rc6�D+�}��8����r���Ɋj&�|����.r>�|:|�Qy�.T|(B�����H�+����R�ΎvM,e`��/qJ�yYB�k�-��ɮ��7(�$� ���CA�<$�>�;?�5ڼ�3�L�b��D*�EZ �U�2?o�<�qϐ�|��~v'�FBR;��fI�4�|I��G��)<-��ံ.`�y o4����F�Wek�^�u	�Zr�k�zO� &��:M~��C�OA�"w�kȽ����a�D�4��ds[�R#&�����6��Iw��3��H(�z˱��a~����f�'i�Qi�ƿg�%/*#�KT�e/�}��<��xbu�x��C�xc�����o���G;�<wH!+?˶>�I@��,+�jK��gv	{���N&�/ 87ze^��}�P��3b���@�������:�k^����
��G-J6u6�)�2��L줟�V�@'��®�D��偨�EqD�k)I��v0�DX�F�Tf~jO��I�E�?r��J�{s ���Y��\�쭺Đ��-+��Jǩ1yS��9%�!�Å��������0s0�gi����ZĖ�0�1�Mxc����1X?��Y���-��f���pS�0
Z�Gui��g�z<�_�L� ��-����N2�p
m�&�F	#�H��}/f�1����B�f�U�C��\��9�HD���m]rk{wIYl��[�O����~O�7{jTb΄��ӌ������;̾Ff5��t�{�M�盉�>�3 �J%|�Ǳ�^�ڲL�t!zt�eK�A��Ϻ�"y�
�>F�ޒEge���V��sf*
ч8&}�7`��S�Yᰫ��X�L+'�����ζ��.J��ZG�$,��
��t�"�P0��[��ٞ�$�J\��+u^�D}nD��a�?��6�"�S�����8{�%�u�N����T���ڎ�b�9�F7�v_S�>7_��:�Nre[�9��
�MLw�l�(�%GݩK�Vu����T�@�j{���[��K}���Y�!����L�<�-�S9��;+N=�������Uc���T�U�4��~b%���PS�`��-)*@��ݲd����a��4�Y����~Lu�1 b�Dw��͒_V��+w�F����-�.�_9Һ�>��?�*.�V���;��7nЫO��+�������+�W�Z��:x����+Xȿ��6�_��L
W��a8�m�퟼uc�-�H��Z���ڐᲃf��"�x+�j(��7Q^�c�@���#:7*�(�`����~��?//#���NX�׈����j��BJ�./7HP���V5�[�j��t��8�e�������HV�n7 X+S�輊!`U쩶� �ðD������"�yaK�e�"C��1 _���&�þ� xg��qf����\�����(�u�Uπ\ ��7�����܆��z��p,0G�%<�۰�GHKĬV�.Oׁא	v�֝���X����D8,)��L����>��Z���>1�Ұ?��8��W��ݚ�����/�����1�����J-��i�|x�[F�l��w4�F�0�`'�C=�d�sF
�A��̣%7�����8��y��f�)I.y��ˇ2Y/>kL��1g�NĬ��*B�1�McdJ֡2��Y�[��D.�K=zT�ٳU�>)��lI��ɞ��ꉜ���y&5k0x�4�#�����S�Z"��D��Ø�I|װ�5�K�PBa���g��0�-%���jn�-�E�=��v�O����6�*:��D��t8CK�r`@MI�iRxkK)�"��!��ʵۭ�:�= m�� 1T��l�Of�Ч��	 &ƥ���6�<@6�gT��ACP�^��Z� �dZ�E�S�c�2�Odĺ�&>C���g�Ѿ���!^�C�s��sd��&���8�ow�������;
�Esae�K��ey�P�1W�QV�ͧk�mG�`N��H��Kȕ����8��ɟ�AS0k�=|5%Eǥ����@�A<0��VM�x%���}�/e��5��_���EQE-ӣwO�'_�ggȌ\8X[�ǅ�ǨS��S�L��Z�v����-O:*���ǯ��i�nC�gV��K����{�p+"��/v���L��]r�A�/+B�,��E�(�~m�F��a�dʷ���@�W�X&D]�%MX�fo!�P�0M���]�`,�a`H�5�rQ�Y{�#soҾ�/V��F)���uW�DҬ�:.T3)ZS�$b�jD�����K�m;%��J�#��$��1N�	������Վ%�)��:	9����F,7g��[�ns������e:AgH˷ ��[�g��L'��SY��wխ���tݙչ �x�|���i6�b�[bȌS�����:��*���S���]c�s��R�u��x[�8{�䤆H�Cv��Y�'��C���G��?dB�d�Gɿ�Ў�oϐ2�����S�\�f���}��Pɹ>�>���p>�/���f��KI4Lvv�6ٛs����W��b*WL�Cwbs�W�/��m��k�G��&ߊ6a���F�������BAX�(�M�U���\���`ϩD�|zM�۸O��2:���I���� �ET�������8�P����|�M�f���x\Q�K�x��f0_E�E;�A�v9�cd�$�z7�x�4�#��+n� �q�H����Vz�?��a�����b�"���9���(*�㕇��o#-x�wZ#����]A��g���&��3r�(Ĳ
SE1���OA{4#3�;�&���ޡ�P��.f�7vb.�fw�34���/u5h�<1)��}��R��n�/ƃ��N؎�2R��~�>g�X��q_""M�	���f7~_k��G��%h��N�8�@g�+j�|�u6��6��E���gt�d%�J����5%	����H�G���:]�Ҩ9�dIWNxK'^5�-��"ȄdѰ<؀q�^�δ�(���+��������r�F%]y�b*���UFe����kP�򷴏LH<JL��*y��z�����Q�'̺�K�]iF������� |P4��)}bb��_ږ��)Ώ��;6�9�3��/�`Vt���ڊMi�����w���mgЩ`m�~��u�QNg�oS�ģA�&ˈ�y�Dٟ����J�����SH������+���� *H��ǀ�`��
+B��j��M�m�7�o�"�{=�cZ�{�7�G��0��pj�������F���i܈�2�V�<	�l�?̸�oH�- ���{�x�`�����~>s���4�x��C{�%�|��M��@��!���Q��Y�(�oGAa�s\&��2�|)�&�qo[fD��{��6�½����d�:���h�y)^�+�Ư�Z�[gzY�ظ�V��pqz�,ݵ����SV�<:�8r*����~�� Xp9z��r�`������kF��I�v.�6��RT�"�s������ʴ72����ɍ�(IB�P��అRZ	��6�0h~ә	��;��v�k.� ~����{o;��G�z��L��Nz�f"o�|���E+\k�����3ȳ���w��,�-^b*�X�=~���M�f�,��K���q��T�.|��r�a76��.8(4(�
�w�'�8h_�Ϲ[�湐�p��4e*E�4�%a=z�+�[�v�������&�،��L"=��g1n=}���,��<c�Ot?����`'Ȇ�e�NJ�aj
p
�@�LI7�������N~,P�s2]�ibE�0����0N�b����~��Ԅ��8k�l�{>@��L�Aq+�n��c�7b���4 uKΩ]�kdQ�h�#}�A�L�4+��;r�H��3-]T0������4� ^=5�������V�CK�X��C#����%-r����ĺ��a�P���b�h� �N7BY��W�}��4I�-KWQ@����Z�-��[�e��O���1��y�7��JT�u�/ X�X}�]�{�vnG[T\F�EM����wc����2Ca5�D;h�zsפoє�Z���[1L�A�z���{L�,���s�6.&0��a��8]m�y�q�`�t#Gb��Յ6�gT��!���ʶ�8�ߡ�IET.�׽Pk�D�F�2���>�vp���9U�M�(���h1S*��r���%��̂~��Zc���e�=>����T�}
��a�d��4W�N|����E���4~����m�Qv���F����?� �VIE,��!���Σ���W���3ZrK�u���d�82d��z<���X���J����E��ZC�f��4���Z]�� V��P����Ҙ����[y6`유4���ޅ_9�,���ʕ`�'��*םXǄd&������*�.R
8�Yf6x3V=h��xE6�m�6�
LI�c43�	�ض��E�4���$NX-T<�b���N�d+�}*��t��y,��8��p'�������&���ZT� -ݱ|,���s���lE�z��&(�@QFۏ_"�IX��H�w2܆M&�/�m��À�fv�	��4q�)P7���%&���$��g�f<�k'9:�����[��-�F^������W��D8�0)7��"����#�ͤ-��=�I��qwv��;�vVS�Q`L���A}�
�B���c-��O�	
���@�,�R����Q��.��y�+T������pLv71�V��|�p>� �t�"�mSx�j�D�2�z$����\��"Tm�N6X�� ��:�{������c�/_�g���8�RhB`cr'<���:b%F󙥔���$�@��!�~��j����F9j��Yd�+��y{`��Z���ZZ#b�0=p	�'�.t�禪�ŗ���h-�7 KC�ú����{�N�)��p��rv�߽������57<�<@Q-�n���q��ܤ�A��`��l-�,���&�J�D��W�[�v�E�:@d5�_�m�h����*%��\�~�z����$��]�a
΁�퉵-��j��u����o"�C�����MLɭ�6�y�|�+�F�+-gRX17��[;P�|�y���<�$�WR���e;{]�㦮�,���c�̏�l^O;m���|� ��1/��g�&��'�h�
���$k��
����0�<[� G���V%�n�<}~���W"��FX
��Wط�{�mnڭ�?h��Z+a D����!��͚������(�ZI{�|���ޅ�јf��m-�ZH6�$^�n����3���xq�Y+S���g�i㖞/��'g3;������(�ocGw�ȅ�K�y�	�?���0��si?��3��R>H9��_��2�h�y<��JЃ�B_�}ZK%���됹�?R���c^����!n�m=d4Űل�|���Ŕ���x)�o��ϻ������t�s��o�߲��QV���L���QO�<O�ԛѝ��x�z;���Ie:�5w��B3Yu�5���p`� k����2�nf�c)�mr=DYݪ;V�[2���#�(�jO��]���R�z��Ќ"w�Md۠m�p��/�?m�$��,[������~�4����V�-BL�B�cC�9W�����
s�,:�p�26�2�4C8 ����ꐚ�%:��P���JL���z�~����j���M��[�s�ט��Zuo<����%�_�71�O���逝,�TX"�\�OZJ�kL�HK@��"D��(�s�Xs�0w��8�cD��� $�� �6�&4h<^���"DϢ-�D��[��O��'�H�VmvI���P�ސ����� _�ӎV��u�����34�6As<c$�s�'����YI��چ.�2���߃fWԶc��]c:�z�,��'`y���y4����l�ب��=Hp��Q����gX<�/0��l���4>�%	�}%�_�gW,��"���g^�;eZ���1%^O�lA�R��}$��?��g���<ʌZ>?�=�x�0�{�x�$6�n0N��Z.k��(�iGj�x�	����)x=�� ��eч"�Э[�}�=�J���{qqb ~g$����f�����L�L<'�P�����N{w_-4m�¸�%g%«i�V��'����%#����OEp7��.N�z�����3_N-��aQ�Z6 {_d���=� ��{�_��CM;Pv9�Q�xA�M7
��D��?[���QM�k C- �����%%7n��S뇉yT7�o/��OO�ĥ�wja��&���t�'5�����Gf�A�#f��=��cj��`G�`եT:'��YD��a���kt���;Ĺ!� ���P&�~�ʺQݡ�b �"1@Ն�$鮿O�ʑ'�b��&����+Oòp���n��?:���@_��Jь�r��"��Ԧ)��ZI3�\/H�do;����S~��G�3�B_�sX
�Jّ�d�fh�[=@fT���cLM{�;v��9���s�}YW>�I,�ea���b,�>�V&m�S?�\�����_ׅ�4s?�]JqF��B�;��2i-xg����o�i���*T9�*�G��]+�+�@�ע�z�K2�R��f�Ý���]/$�6u �X`����l��S�!����.U� �Oh��6cl 8���+�ө�a����NI��/�Vj������o)3��*�}�y��'Zd��N"T�Od̑��	�E�kJ#�7Ec���(�����A��B�?��Weɺ�E��,��,�{f�s�C#My�"p@A��7w�[�t�(��nH���!-q�E��V���3C�I)�(�qS�A�YF��,�_���_s4̵��~�{�l��3C���k5*VsuA���Mʞ6��V�vH�K~�r��hwr�4��٭������P�]����X�i��!�l�k�Y����f�o�E�Y�X��S0�N�3�Qf��
f��k�7�}�B��^ӆ
�����S�08զ$v�W��2@'k/���n�|��BPӳ%�X��S�,x580.���4���v�T�n�M�@
f߮�;ȫ�'s��v,Q~:ϲ�y�6���u##L��e!?�yy��K�����3�A�_�����
y3��6�2�ϡ�8��|�O��&����JB����;�CS6�U���k�Ho蜧0�� �)�8������F��S��W�LaP��ki%+>�0�i����Rf�{�x���;"@��驕��m �K��e���(4�;���7�b̂Z0bQ�i�tɶ��|�<��Zl�WKǮf-J=�u���C��SlpY����:�R�n���ɋDB@ւ�q
|G���%<FiyEw5W�%N�[ZW�Z� ����}�f�h�����|���$���ɓ|^�أB�+��9�"���b43���*�7���R��u�BG$��"����f&��6]�����_����L�1臰�����A�L��|C��Y��hZ�����1)�)�wbp
���)Q��GX۵n�{��y��Z�
��&ߑޖq��z��J�}V[c2�X��I��w�Ra���زMu���d*l�����$(�3E���I�^�����B�tb�u�$��_�`xq��u��%=KX�R��4�]�ݷ�h�V��W�\S��B�@�ӵ`=��x܎Qs%N�e���|�'���
ek���B-@�g`�5�ziWP�=��<�c����u�kA@��>��Hj�}���gÎ�%�
fR`3 ���vO<tq+�jҍ���+8/Q����y�r|. �'-���0��b�!��.��5��4q"E�N6;/�S��&���-2�]���[0��v��	]!��ru�V��WXgm8Q§�'��G���ˢ�IT	=<n�>����Gg�/�6_,4��kB�H��~eG���:�֠�U��1ɑ��H^��)̌�5#W�kPr�t��"Tw����G믓c�^P�\Ί�3��N�R�<�d�8ǹ״)a���cq�h��b�&<n�ǘ��2���,��{ӛ�kՠ+N@�O�U�_aB���ְW�����X�{���o��YO(|o&����#�+�jT�=�Ik�~7v�W!��Jp��\�-.��n�B=Y!v�C��%�4/�,��Gbu!��LV p��B*��U�	���� ��d�A�,���7@��Io�D)�ӌm��ε��m��A)�.��
z�D��dC*!9�L�� �����5!�=dϺ		��&�W���x�@CņJ]�O�}ԚK;L)�?�������k1�9
�q6C��;��4}i\1�x{ �* w�.�r1o�;7Y�����C7	�� ���Ow�[���?�b5����흽�����]n���<�0va7單��I��R1��]0����K+�Mo���
�<Es�E�2�F/��}3NP�$;�-m{�r��_��?d����"�Ήn���ͣ9<�{E���_�%s:�#�d���}�{x����a���P��U#�3.���ZH����zi����ܧ��򜏃��Y�&��ne�J-W�y�T�i�+~�	X�]���h`O�ybZ|����Tr��J�X�(�3�d�9��'��� ��=����4�&J�Ç��nU%٢�}�z�L�e�c�H\��8�t�b�?�ކ�FG� ~'y�o�B��C������4��[�*8�B"	N��"0���Sa� ����w�oy�R{�k=۫䴹�2���Fm�ǆ7�0x|͉X@�Vy����0��UA�3�yݻ络�ݜ+�Mc���T�?�[��g��v��T6bw\��� XY����V�p��ȡ%��]e:SE��\E�B��0��R���H�]4� �0_�dz@�̌�k��#.w��M6�콩��!���p�$��1���j�Mp���,C�`�� O�ɭ��,C��S���2x*���ցR?C�9�;~��>�h��M~�(��g�_^����:���d|R19߈�QhK��Q/ٍW��#D�w@uJ��?��$��e�:����`ƀ�7�J�s(Tw�?VdR �ӪVG���]`!P�<&�!�ܼզn�1 �a�5(�1��~�Q4��?4�
eV�N{Q�jR���!9��Cǖgu��mG��~��75N��Tgv�@tl�8�k����s8~ʊ�|Vv��ل$^�#�Φ*獜�T������T��)~�h�}첾*����j�C�8L���k�˔!ϔ&E���PW��T]u{wK��~`&!�:hh�� �a`�S�nAȪ��'���u���BK`;�d�TJ�������>��10�1�4s�'�*�-S�s��J�I�����oec>���P�\�Uz�a}!n�Z�M�о�(�x\T3&�\��mg2�R#<�!5�	���W ��{��.���D���Q���<;;��o����v�/@�(p�My���pw�	5=��p|zk��F��%�m�ܤ*����!;�$_��}�-ّs+Sn�ǐ�����$dXCY^�����[��J�`"���aѽ� iAY�YH��-WA�M?��{_/��Ẍ́�}�݀���8�3�؎̕��mg˪�k�,���h��j�-���OY^��]�ߡ
���ΔK�e:P�m��KV�9�s�x�|�Q|���.:�bI ��D���W1j�=�}4	���(f("��FA8V�v��G֛0���Y��?�А�S%m<������f�
��G��������O),p�f���S���JV0����h�^�mZ�_��`i>Z�҃y���[�uI�c���Us�e��腗�d4n��xv~'���Fr�u.��
9Yh3Rl�q�������B6��&º�e�m�bp�eot�ЩEHt@Wi�
_�҂>0[\L[;�+���+�Ԇܜ3i�=~��7�6?͊�j��˷�7ce����JϪ��k	���_TT�<��+���8�=�8��%��T�Y�5���Gn]^1d���_q����32= ^a�e�Ģ�+���w�lH�I��8@��5��t�)|� X��T�����12;�P��T�+d�7�\%�����?)]żX��&�����Aƃݯ�Rj�l�1��v�Є����?�W?w;�2(��jj�����q�/����V�����SY���f]��UY��r�8\��P��*N	Aɉ�^<Sl0~Y�N�ʋ[�*s����Ex���d��'��.B4�7An��uL.F�o���7(Px;���ׁ�b�g�J���8�by��t��rYH=��=�J�U���������%'ۤ����t�l�{��h�(T�Qw�G��D&��*e�Jl+s���v
I>�"��*ԈVt!�Nj�՛���:�.r&��v|m���[�ԃ����&���*ѥ�	�Ki�ݻJ̨398Q�ދ*FI���v	���	�Z*��r�=��N(�t�C���ZB~C0���Z-�����+��X��\�G��NX�s/=(z��nV,��aϴt�_�N��V�]@�ȩ����v�5~bL�����N=��D�G��X�̣�O�����Za������dUfF�y��$��H(�蚨�	h뽏�-��.����<�����}_�7o羏�)���z��b=�G��4�8�&��:��1xĂ����Bdl����#�`�Z���`W�Ty|J��6K���Dv��mͰ-J��vy[y5X�sI��4�R%@�~��Yn�v��t;�P�ZzPA|Q���@,�{���31�*aD�C���mˇ�c��<��J�G{u�T�hgs����m����g��T�R��[.V��ow��x�b.���Y��5*���vZ�UO�K�PB~����;x)>��MUJY� �m��7)�}D��O�@���aW6.baֲ�~�ǷT��FBۿ���5�T-�y�M�RT��Q��X~c�i6� ���T��I�)��xB9g4Tf����QX�����oj����� 	@�Y��bX�4��A����e}��.��q �]�+-$_��I3Ie�cVr�n �h�-�sCC,�*����v��܎���A6M�M#�jp��O��F�d�QaB��"��R�/�!Wшz��d󵓌~�>��+F��mV8�K��/f�,K�>c�}�d�5E���p$K"_Z(�U�a��lA�1]q�h%��Մ�ȔѦ��y��D�O�{w��7�1(!���e!d�� �q��j��@D����cy%���|s��N�"QF;Z�+l%��"�= �')�C8�<A
0�򫲡ϬT�J}�õ�l����;���okڒ�V�\#b��>� �R����Q�q�����$$�\!��)�~���#.DoRs]���e/���
b`*��?J�°ogK�`�tw�CL�%�%D�DCG�ק���Be�:������LRtGaL��?�8^�<U�����@J1����%��T���Z�'������d�/.f^Y}%�G�Z��74���1���*��.=���Ow�ͩ�7��n>����_�ͤt��#�m�[9�f����Q�㲕:���WO�y���^N�-���P)�� q=�zD�7a>R%�}6�ٙ��WȻ�[6(I�e��j+4����Z�w�N��M�+��?��d@W��UD��D�c.�����W|o�e�h�E!*U�=Xkg'�����r�z:�S��Un[-k��{L3=�����|�7����rm�@k��w���܇GٵvΕ�<�0szjD���B�Vav4pTX���_p��3�sj�;����G��@@���(��I;I`-%7"@_�3��)%�1�.��$a�ꉻ�G�,Q�(^՝+�*����_{K��~:��ˇX��i�Nz���Z�8`*���L�)��������!���H ]J%�k��t~в���z��0Vى漘`VQ�D��W-�s������f��i3oN�Ѭ�à0(��CBU����Q�Qբ�2q���GF�����-��>{�D�i[�z�"���X��:�����y��͓���zn�g�����$���}w��yo$�u���U��T�)T#ɀs�`�Xj�?�l�lF%�"��C������bC#i�
t�R��,����J�6�yLa1�# Q�[Y����|��:�����19n���sZ�vЈ��o��}�5}(Ejx6C/���Ar���<�C�P!7��3�N��*}鵆j���Ͷ��ý�Ò�=�3i��
h�^ #qVJx�hf7;��b���)ӟU�5�E<S=~*���n#�`|��xZ���0��|�Ť�G�Lǒ���6����5u���Q!�B�ޚ����%-3(����b���D])�����v�7���X���L��@!�d����q��+��sz2-m�!GGO໮�"�P,�1d�H���o�'���!����J),j͹d �
�mI���%żK�C+逧
�3�f���z��$��A���ĺ��[<��ԧ/�����^ҕ�s�s@�oŻq;�����Y��X��j_�L���g�E⼨,͇H�	˾�6YE[��r��{,ʶ��> `�����K�Ã�/�(�/�º2��-��I�6LGq��>G8�hHQ�kƹ�+�6L�A�m"Toey�\�Jf���y�x7��fyɻN��6V��l���W^�����e�����hy��OR�⋜Dl��:��x���~�V��(�ʊyi���},
wob��j��<m�_�#V5<��O��/��}e��0c�ܮ��IG�8��w�I#@
+n�/�N�j�O,�*\s��hnv�ⱃ�e����z�cLկ��sd�n�WCH}��2^׋�U[��i9V�;��5�X����#�/ɻbH����P�TM͂��8}�IČ�;\�*�dי��L�]��E�6y,2����q/�OQ�G�;r�Ok�m��=AԖ���:t1-	9,� ���S F^� nе��'Mvc:��e�􆞚�=@�8�4I2��*_/��.T�����&Y6��>=
��#8j�⇗غO�����"�G&	�96cq*���ЬZ��7�2�H��*�
��2������@4��C�PH� o�O@8��������_�l�n/���߁G�O9��Ҟͦ`IY�3�y�6T�_������J���7᜖�N��dL���Et&*�?���mе���Eq���z*��81y�/����M�]�ϯ� �ʉ��8��� �;�^���+�+��a���:�pl�
m�1x���E����ř���dkZ��ǡzZQԅa؈�<NgC���eu46}:��`k��kM�D �k�x���j�&;����t ������!�q�VDA�f3�b�迒�ٍn1���[h`qkPB�A{��벘�{�a�>N�)�y��+F�{c�n���w��r��79��J�V(�zm�O&=�Պ��A͎��$y 
9�ց&�V(@�+�����@̛����r"6�Yi�������L7*cK	F<!G����8�ѪW F�.ATJp���ϳ�аs���Ͻ:ݺy\{eo&$>�L�{��
.��5�ς��%��*"o���ge"��U0d:k�؝i\N�ۈ�ޞ�Ω���� ����-
2����cר6����Fɠ�ә����ZLL����9� �����v��z�b�y��]�jW,Dy���D�a����f��\�w��my�����%� p<<�̀�����5;1ь�Q;����[#=��g�{�pC�i��,���ɷU�T��b���6����7om|����I}��G���_Ŀ��Q9���d���|^
e�{疱��m0\�b:�e��݀]�l�Ţ=�D�E�҇H$�濭���2����7=�K�aYu�b��τS�g9�/D���~3�������qaz�R��A$� ����@劍��.��㘊=�N\MCrw�T¤��|#�mB�����0�u�|D�`3�n4�4
���/�ٸH�XA<'  =.�4>�;�Rk6oI�p���gc������[aׁ`��1g�]),5�?�m'H��r��>�++@_+Ŝ���)�7�c��>ۥ�_M:{n�2����S:i�[�F�_dV�"os�{J�g�1=��8�]�<[��(4ӽ���<9���I�DEh���j�Nr,:Q*�c(���G�y[�w?��}ZT�ކ�j1��/�����0Ml@��c��kWqk:�b�pL�r��}6���+��5���M��׈/�EO��w�Yz�Xh��=���2����{?�~@����H1���dD ��,�I��w�U�2�E����q�:ux`���"�a����,ͅ&t�n���p�)Z��Df�2n�?���C��YE�/$��=w#C~�N�[�J�����zõ, �}Bǣ�[�@�����:�T�5W��W��O4� ��1T������|�B��y�ah ω���M�t0l�W��_��Ai	���[��ϒ����-�X(P��S������z蚛�"���)@��M]���Eߙ8��ҁ{5[|��U-�I��=Ne�ɋ�x�i-�y[�7>�K�$��E�\�p2PRQ)���h�M�����d�ø(-�"e���]��-���������=ȥ��C`��\�J�j���Ar6�T�_���������74���v�+[B1�Pg	��\F�F��A��������3����m��`j�Ѳ��8��Bݨ��|���J�^�)L�$\���T�PIJ��	�fK��.�>�9���.�C6ӮW��p�-����j��HSL�>������ip�:�i R}��9{'jͯ[f/f�H�"Nd���V�Y��n��Գ�pc �J�r����p�m�<�5�:'��V��or\�p�u���s���I$�a���6�.�S(�y:�ME ��� ��̠DH�z���ڰ¶~�jc^#���$��@J^�4/� 	�����I�X��uH���r�g�
�:oË���H_��I�J�AD����*2
�a��ٶq���-)�4;�pw��m��B��Dr���V6��1���f�'@����4=�����mӿ0���BZ����-+b̸J�����o׺�lx����E��Qϒ��8Y>�����*�m�1H�sp��u5>��k{����$�/n ����D�>c��s�SW��E�:� \|U�J� ���M�m�fb��Q��m�[N��B�Jk�Y��=dd��D޷�4V
��C�x�`��&���^B�-�qVR��k�Z��M��=��mWQdHoOH�F�mSD�ͦs���]���\�Ѝtz��\y*��Ѣr{���U��.��AN�OH�Q��b����J�414b����f�5R��U����fm����3��E<{���[s|QܣȔ"���Qjʱ��w����t�ٚ��e.�~I�fg^�ܒI�57�Z��U�!96�o�7�Y��b�:��h�"wR�+���k�@�[�柔��>_�y������Ms���T�����?Q4�s�&;Y�H�q�@�כ:0ف�����#��f����cm9ge�xi�-���R����Z��Sz�N[P(���uz(la[!�L�~\fg��B3���v����e�O�i��� J�w��/��BFL�iA�Hk5h""b�b�=M~�o�

S�Fq3�Rŋ�!���0�D�WԠ(#�{��/kΥ5:QùF��4��| �ڡV�k�=����(��2k���S�8\��w�����k��qO�KZ؁O�Vg�ܷi��:k������t5�lA�;Kn~A��`�0ĕg����d����&NQG
Hi���4?�v0\���n��^�$bl�	<�K>5��mz�"�[�� ��)@.l���:�C�q�hOH'�� ���Iǀ��Sy_C��� JU�A�#6�Xm��;�s���,t�{3r�W�8h�_�O�~s�P�!)�0NM ����Y�nv'y,� Y��s�����k	|�CR�A��0�]'�k�J�$�Z��L������K�X��a"]D>�S}�J>}�����?N��A�wѤ�3K>�(à�W�i��U
�5����C+��GP{�!�y�����$/�̂����vԸ���v�;�G��zRI7MlaC\�:�]�`f��S)� �ґo*di7띮ģ�ﻺ�si!����/�)[��R��sȄ��&T�)�i��^�ɴ�RQ�<Dw���j#��g���z~�f@��?�&��[�U	G$��":D����m�+�s&s�u�Z�/�]тR��3<���?5���B�dW��-�I�]&}�����:�ܴ?�d<읊#�-�p�Z"ME�F�i�9�R�=1u���=�"�ZQ��]��Iؠ/"nB᳙9j�Sf*�ٱ8����C��/t%r�h��Ҧs����|*}<�
R@�q���sQd!)�g��^���p0}3o._�<?>`d^K����+�Z1�e8��3��F셄�r�(ڊx�,����	�	�L��,�j�Jn�S���A_t���'	u�Հ�5ѿ�B]lP���?`��MU$���$Po��?z�|h���[�L~���^X�r��=F��0ϸ4F��JX�~X��X�K�����������7�ށ���ؘ�="���#_U!����*&H�D/��#���A*��-��et�
o�&3F�&8IB{f��������0���9G���h�;�? �[�u�m��C�����0UW4SPdE��y�W�jI�sXOU �+
P4��~a!��b�o��P�Dt���t�4�����d��s�%q>�����GPt0�.�NW4$���:9�,��[�lP���D��h��*4��d�����@�	��g=�4�2���Z7(莽ש����}�mw(���y�tr偁�j�f��E+�q�8�!��^�}�yAg�.��-���Sd���.����Ӎ���)]d�Q������3�f��U�*�9-�"tg�C��Lm��6����c�J2�FD��]�M`�ͽ�P�S2`e��M.B ������m���ռ�=w�t�3��گ�5��rO��Q���/"�]����E�v��( rx�R�<��UMY_�Y�QCV�1O���7�v`�=�F��
v�Y�A��v���D�g��&�RE��E����4m>����a}��'����Ѩ�eu`F��*%�W�5�eF��[vŗ���� ��K�mV����Ң_])��{1�;�.�2Bu�G�P4ᔬ`�.Y8��I��ef|�_t4�+�#L��t�3���k*��)���li�^�6CM�F;^9Sߡ�� 8
�Z�^o�h�k`�g��a��ȍzK��S���t��P��H?Ἀ'.�v�na��E���o�>S�	�*�<S�0�&C��l� ܂6f��VD���.��o��&f�����D�p	�}^ᥭC���&��`6��Y��*�'B���ȱyZ�YZ���$���)�W�Ϗ�7��qt�hV#�"��u���w���S��M�����ۙK���ɏ)�U�P�VV�����M�(���ee�ǖ�8����eo��f,	�E�h��c'���g�O��w������H����Ɇ�c�0�!� :�J�x�|n/��jk+�afx��[kW�R����Ѥ�Ώ��_���2)��sŁ�O���W�'��W��rQ�?�$���@��"U�q�����S/: ,���/�K��!a:W��Ea�n�>�%.雅ۀ���^�ɟv2��]m���l�����w�sG����Ȱ��l�;�B�$��[�F��R��s2�0Y�엻U���W���c&�A3�߲_8���S����{�>n4hL"�M�I|,�{���9|D�]��q�Z*�1���V-�WZ]��N�9�\�J�I�mm����s������T�(���J�5����"i���^�^�qk�����z������,���L��]�bRL���T%� _�՗N�7�����`�b�?���'A��ۍ�l��ǆD�| ����A�]���>�MO��XS�vw�\���HF��ڎ_4�5��ޖ�xl{��V1��)��=�!��t^�a1;���z ��O2���<ӷk�肾��??x�h��m�K�<�_���bTJR|�ׅ�I�I{�*x-��L��l���E���N;����Nm2Nh��λ H����f?��P�
3����E)?V:<ș��r�ާ�BI[��~ikD95�H�VO�n����	��0�s�љ�-�1�G
Y�VV%�M��c���������'�����8!�.>bp��Y�	��=�bzj� 6mJ��� ~7��Y�n[n;�H~rg|&7�`��ik&�lX�G�����f��سeA�CE\8���N�v����o��Gz�N�^�E�����+wf�)b�L��~կ4z~%����@u��o��sSs:��.ߊƺz��h|����DQ��j">[J!�Yl�BU��֞K&܃Yw�<��,2�s�밿K�*��e�v~I�)/��?ծ����`+/�b+q�ahB��a ���R�9c�_*�X%���_�X��B�*��[��H��ĴM�{��}Uz~$�C<;�&+�����r`"�zɈ�N�0��,]ry$9�'��F�8Uۓ�	/܄� �e/_B!}ͪ'sr`��q G�>4X�)�0�8��B�@W�/$y�X!Ɓ�� K��g��˅��p\��0i���}�sA 	Rw.�K�⻪D=s]�����~�3�Q^@ �9jwy�ߧ$�k�_c�c�5�;-�qA���}W!��)�V��y�^駨�����SuQ̾dŶ+;�.,�(ڂ�T��6@��Q*�Q����y�uX���d
e��`�92f
�&D76\�8��\sq"w�ަD�YL�qJ+~0z�-)u9���7&���y�Mx �u��ёT���|x��:�C7���J�zY�x��u��/�"�cP�� �iC7�$;z�[��F�<
/�ҏ+�� �f�>n���|]{t(�L�-�rt���J��wR0���+��;�����ń�|����L&�@>S&G���ez�y�@�1B�M12�i�\���=$�p<�oIL��xw�j�a�T�jX���h�Q�4��9j��{YV�dث�9G׹��aǦdڠ��W��(3�t���NdW�f^��.���~��Rf-�IXl,v�3ٱ��`��+�e�뀩�Z&B�#��yA���Ɲ����Q���	�Ԫ̏��G�� e��9�7��"������]w�i��}��+Φ�}���[����5�o(�@+�k��T|��2�`!�oח��;��J�`w����~&	�k<�Q�g�X���ݬ����[�H1&�p3O x�����6ŴG}�XP��S�@����S�Ϭ5��"�*ہ^Ӳ,�e�9 �Ac�BI�
��w����a_�lNb/�p&]��d �be�p�.��@5%p��d�������́��'�+ʥg�\e
"��|�8�� ��·��`��)6�@I?��p��پ�fX=z���SYYw;��!2�%�m�����lFY���q��g�w�>!�i�/���������H������̉��@���/�0�S+<���D��~�`9�*�+ry�N�b-e3�j��dw���x4v�g(����`�u>�c�L
�1j׫1֧�#}r���_���w{��jp����0�ˇ��>�&����<��n�4���RI�l?���4#ړm! )�)/f�#׳	�	�y��� :��\���,�GY�G-�mYQ�@E�P��&"�WO�/<�Ȧ:�����fy�Yp�� |u>�G��i!2���BS7���R������6���s9�ze�h[�{�y��^\�W���ݲgWA%��)�u���W�q��9�r�n��f��C�_���
�zE����j�կ�D_,AX������MGj�!��ɮV�^e���"�Yk1�/��D�E�p��S�6~y�b>����O��9.z���MW	h"k��Z%C�#"Qu�rǮ}NK���l���$	3X�)u�������oB��+LT�ŇK�!��H���L��������aQqX�����B%�+�����{+��䡆=B�}0%GE��P�����_H���F��p߃�%���:�&<�-ٮ\B"$߇ܘx Q����3�/eo	�	����� '����}�B�;�"��z)�H�7".���wO�r�e|��`7���W��jd�:}MD+�a��Ъ��{ ]�iî=��*��Ac�j�ל=[	����������ö ��b�x�҃Y�l�S"�\�5�1ǛA�ޒ�J98�q[����&EМ=�2C;�6�dj'�D0Է�/בD�O��/$�?�Z��j��EXM�'�?!acm�]v41"���#>.��2���MU+�<��L+��w��zİ�sK�u?�B?�w���5���hrٝ��]����wb���J�sp�ܒ���v��0X2�	]j��2C��2�@�	Tw�A��ҾJ��jQt�[�~g�Xa+�?�8�"�(���$���D�`��7ڭ>��8	V�_��;w��`p1��(�0���`y��ˁ��	�r5��γ@�+����D8;������1*n���4����g��"߸ň���C��s���}f�;�GZ� �թҘ��s�]ëK�19{_<��rF3�R=]�W��	0�v~h�8�H�G޸l�gxKF|8�ZP[g7@A���~�S�۳��Ɋ��"�Z,�m�sL��f��I�7>�I��K�cH�Sv%�u��Q�&�(�]]����u��\�Oإ��X�vxd��� �T��=0������	�r�-�x�ԌTz�X�� �-eyg;�Hw�}Eo���QrS�9h��������b�v��r[��o�: ���%�b^=~_�uA��ȸ��O�sW��I�l�o�X Y���P�,`��0~�٩��"�|���T֠f��L�w�I�V�tx4�a*O��SȷaFB����`��2���t��8�˸Cp�;���)��G�u��8��Zr�M�]@�A���I,�ջ��BNS �U�zD��ZX<uA���:k��,֒�Ҿ	�������������q-�O���x�ɓ��`�"�Ӏ��b����_���>D��G�ͷ;�XJ-�?�~b%��%`GN�y�8ˌ�Tk
5�����>�1������pz ��+B��
���#?��6H��X.��bg����_��ZXZ.UPX���S
@o���=�'xt ��n�hl�(� 8��*�"��I)�	��k\a������$x/{Ž��y��%u|��k�*b#k3��� n��{^8ݨ�`�g�fUv�(b՝��rU_�{vC���ĵݡ�U����t��Y�W^(w���7��g�_^�d��.����3�0�n�o�;z�(P03�M���<���*GO3<�Y�x��kU:�hB6w����p�v�q9��[�����7.H��y��{o_v]D|whK`~㌆��2��Q��I5��:��fYp�i����1��~/���dM����+��myH�2�p�O�8�t�2~WT*�3�=�t�q�7ZP`6H4��2���R�D+��?Ƥ��q7���ɢ�/oBX���O���Gu�'P�m�Z�Os��|>���b���ApԷ���?��H�Cǖ��-���x�$ **�eo����- ),<ɐ�4�G�̎(�����J�����d��gD=y���"ǚ������&I��@B���l`�Y����T�g���Ě���o�J�ޭk�&�i;?���9�b�p4�Bt�L�CJ:��Tl=���/eA����.�M�'��ؽB���O��%�1�sڨ��
OD����"0ܿ��,��qxh��=��-�d(��Y1v���l�o������-A&�ֳT��O9�;I������<����QU)wx��������l�t���E�ϏW֗���T���j8w#��R��')�F�ZȨ���i�ўH�]?�I��۩B���ྜྷ';��?�K�⩑�d	ZJ�j��T�UmX"�a*+)��0z��'¹�}8N���Ҋj`����R8�`F�Rx�[b,�ɂv_��P��aO�R���w��\"K�>ڱ�R]F�'�]��	-�[1�����R���V*���i�'���ly��WA�֊"�q��H�w�����$ ��K���+B�l {6j#����-*B4ɩj �b�nL�u��YQ� N���]Y�Va!!a
R�K�6���x�}
t1B��M'ǩ���v�O�4��13���dQQn����i�����m�~��r�z*���!DTܧ.�oFN�&$%��`�#���pb����h� @tduR_�J�O������+��V���>����۪y��n	Y�D�k��T�~�6�FlU"���7�]�&�y;��kH,��4�á�L��n�&$`�r�wn��I���H�&��]�(��$�- ���^n�������S���
����W��EIu�a���DI��Y�q�7��[3��M�8��ߟf����S��
[Iͭ�}04s�5M{&��Gī�B� N�8�ͺH
V����͞�R��N�@I��0�k�8��e!4 7F4RK���S�KV��G�1 $�B�B4��v�S�&u���)�Ac���M�<d%��KAu����Z���^eeBn��� ���������w>0��)�i�I��Oh6��L�#��yd����>w��S�um7�Z��6�	R�ج
� zdNK�$�����jX= QN¡�3-�J��л9[���?�=4�,�b�b��<7ne��v���)��Y����jZ5���>�@9��b��حQ���!ѫ����.��"�o�\�6u���ۖ��?r2L�"��Em�KT��IcAr�Dl؉����k��}.ӥ����UL�c��� K��lΚ���F�ǽQ��+��_� ��}BT2� ���/pY�s���3���x�'0K�\�)@f�<dzF� Z��a%�Xc�xi����87�wOh���90�� �KAp��ߟ��8#����7��SSQD�n%�� �}_�?si�d4�q�å�O�M���m%����1�@�Z$6���V�Trr͓�� E����'�g�.\>�=%*�O��a��T�eiA��-�~S�Ð=�x⢻|R�9#;��A+6Ś���1��:�B�bQg�A�rѺov\pЌYem���2��z/�|}c҄���I�Z�[��E��l�2V��"P��de"�(%����A'���|A���/��\�p�f8{��):Rj��:��Z�;=I;"��c�8Hf܄A>���ׂ�a��7��r,��Q�i�"�Nc}U�[�M�����O�<� O~�3�Xń��d���K�Xҟ)�� !��z̡�eAs���c��Uk<�l�p�:�%h�e��_Ķ�:-��X�7�w�7�(ҿ������c���Ҝl�>N������3��(%�u%��gu��c�ƷԬ��1�=�7?^�L��
�|��%���[�I��>U�d��8�Ώ2��c��+������%8̓ �Y�+UO�y~W] �+�MF�ż�G����QʼO��V3�$�']��*s	��b:�	JHm�L~VY �8+����rY,,a`�%�o7��3��ω��a<��ʊ�aZc	�m��tK�厕�����ׄ/D�-]�U�
8��X���D��q����h�����S"l��nTs'��}C�QG�4lT��M��m�S�a �����
��%��'����u�r�g���8|�Ͳ������a��9+,����k,�]r?}�t������j�F2�yp,��K1�Ѱ���9�l'���\XG<�����}D��c�T<?m�֤�p �X��ĉ	�0.����.�Yrm�]R�s6mhpz�΃K�����{E6���S���F���=���e[(4Dz�C�M'(g ����Elj����Ī �<���R������������f�>���a���nG88+�UӚ�t��� ���<D�s 7�"������O)�A'�4a�C��ۨ�T��MPz%I��H��Nq����ƒ��+j�3  �<�GwO��gb�&�� >f���se^��9��X|h��S���}
�X�=?�әR�`!�'�X������$�!O3�ރhJx�:H���L�"���Ģ�T�?Q�P�ԍ|��
�Q��;K�k
I��:]g�6�s�s��(�	��`�Sa�ib��7�H<Y�,(މ� ��K3f��m�[�y>_v���CS��Nd_AL(�m/����t���t�s�qhW�f��1���OMԈ�cA��ZCw(���7v>n3��Y4wV�����*����Ƕ���R>�'�I�أ)R��gA�uDM�k���)n�R?>��N��:���F�)�E^<�
	�/$�O�QRW�bH�L���xό�¿�%e���m]���b�^��dq&���Tz���(����T��wR>�Z�i��1s$Ȫǹ;���̏W"A������ K�T ;�m�g����ri���~��9R��$���L��������@��-Ǽ�"�^S��^�f�k��0Sw�S��
\�ɛ��Q�8lʄE�5�FƄ?��a\�� 4��5�Rrw.ȹ��ҾNA�i����ݥ5�C��G��I�-�Մk���;8�o�N��G�9+]���&)x�����ʗ��)�tO-����2$cH��M�Q������Y5�R�I̻\��ښP��� �A�:���M�;����o�Z���Y��^윹kV��ЬU�anz&�~��t���B�[��j����M������ ���E%�������'���\7	:��E�I���!׉���NP�aY�����{|ukTO��bV�Z
o�7��w��y�R���5SC�6�-��kㅸ��B��2"+R����G�`b��ld�L���7x�o$�!64��c�Q�����>r�=o�ǖ���~x�/Jf����}���q�@Z7<-�ꥧ�{�9=DߝW����E|2��=����e�1�g#�$b3U�LN�;��p�	h��Rqd!	��x��"���&^��4�;߮@�ah���"4��j֧����Н�]����x�ʜ�˒Ե1�L�[�RG���(�9wi��c�:�,
2�{��wD�a:��^ovn�������Jְ��A�6O�C��|ɗm������ om���4� �̟�����ɋ��f�~�(�?�ܖ`#xvz������ȕD��9��׻/ײ�N�c�{����:�Ŗb	q;X=�	���3 P�!|9�������-&/��ϟ�)}�wj/�&?DX�7�s_�I�����(<�5ZL�K}C���OQn�{��)bݒ�S����0I�!��]wF_!�m�
9N��a-�05.��Ɖ��#��H�҅�^P��_Ē�<T��%V���H�bh%���e��m�k/}`TN�:�Ԁ��1d�z�D�-lE�]z#�9��>�ᣋ��+#j����v�t��n���]�M�AnEJV��e�Mk��H�@�]��83^o;WQ��(�u�������t��̿$O�������S��	M���h���vy��?W�&AX���f�s~�l �ϔ4��Nv�D�Ω[����{����������y`e�Bk�U��8r�Ĳ��� �i<6�1����g�j�z���A�&����d{�z	��-�Y�,ϟ��y�Eɣ-�W��E[�D��ҫR6�A"�$�m*5e����=/ڒ������������.ܸ�@r7���Bq�u:.Ќ@�,�;~��K�lGkfv1�pj���XS��ꮪ�Yؐs�_::��ϧy9SE������bj����%�I�T3b٩���#�k�����r�Xi���s]5:�il,$=T 6Ĺ�U��x_r<����X�!v�03ݥƃVʨ��L�����Q��i�T(��T�^`�N
ab =n�o�e��ڜY��dW�1��h�����c����7z<I9n��{���ûp��yq����ۭ���0�����<�B��-�_<���`�_�`D\���H�=%l]`|�GZCG #�R h��Z�ڐ�	���'M�(��(]_�=��d+��M���=6�u����XE���d�� 8��f��ȁ�.���XeQ�o	E�3|�O�r�	u���L�n����x���q5�\�=A:��R.�K�P����t��6o���(E�i32��<��C�w0M��I�h؊�9�U���18�%z�p����
f���|~8��s�B�-���¦"��o3N����V紝� �����|O��YbBVm�T��� ��Юş'tT�X+Zk�ڇ)\i,�K&����]����.�����`zǙaQ�S��K�X���mZ�HD�  ��K�x����Q�:p]:ÆVCk�ԯ0��~��'8U��f�s�G`ӎl�p�3Y�D�]�}c7��WKe�][[�E���\;�l~r4���5\�����/�	����$�JHX䛭Wd'ǞI�G�/>��sꞔ-�nP%��Y��G ������a�T2E=�"�pwq�Kf�G��� h�,r^Mn0���3 ��㲮l���]ͤy��$�->WP�gE:z�JWCO#����\�KKD�X8x\N=-�Wpm�>ٕ�Q���£�Fʃ�~(�Z���ӡ�	�d���$�3��&T��pl�QJ����R��-�h$�@���۠�LD���cy �Ё5���qw�1�Z�L�w���0�d�;�{�]�����m��Y�qF�Jf��)����f^�����������{o/+�o4'=�훸D�[��Y[�H`oR�[��b5��s"�[g���-�i��s�Z�?�[s��;=�˿и���C{� .x0ٔ�'�=���5f����Ƹ�Z������7Fl����;��k�I ��9�_魣c�a�߷�#ī��.Փ��\#�@P���f��&�ٲ�K��J�=����}2�}����lK��w�.#��JD�!V[�?�~:]��� .Ν�֪�"��Ek�6yz�2��eͦ<��쭤Q%gc��.u��� o��̈��w�"�p�Ϲڟ��B>$|��k��ы߅��#	�����S�8�\l���n�
�/E��š*?In�2��[�4Ml� n7�+���1�i3�\1�5Ť�IO�.�78��I��� E+�U��.<i�~���u��6/HB:L���x.u�'
y+�6�ĳ��1��b�<����୬��̶ ���]���sv0�lU�	���
��V���c��輹h嘠���~0YidIb�ħ�#e������@�f�UB��i���XH�.�-k��K��RW�x����z����."趏ژrjL(�s�)`����|�?�#uf�d��5�R�Ǫ�a�V���M4X��}j�z2A�S�	�ѻ5�&W2�Ʌqg�Z����m�i���L;�P�M��N׮P�/@�7e+�|F'O�P�f�CV�}Ʌ*���t�CV$g�u.��=�vGNRG��/sX	[YS���
�Ix>`M��PRT��h~�@@`�JPڄ���įu��Z������10b-h�AIJO���V�{�MsڄMs �0��o��蹻��b.��e�ԕ\�7�� T��ywO�+��=&8���i�-; ��ֵ��^����mw�)�*�ZtQ�E
�򭅄�a�Y��2d�K���I8�eC��ߒ��W�5���6���vq��0�&�F�h�#�����~�ZPn��Z���w���܉��i�˨��=#�0��M�I[�rߘ �-#�1]�{_"�rqVMK�;�Vh)0�S������YF��2�G _�S��9���~L�{�v�fa64��&��[��������W�$������%��2�k��qU�ZSH߄�@p�V��s��{m�m�uq3aR���]_���wJҪ5�=EL�B׊D�*��j*�D����p#�WaE�2Oߗգ�P3>x���Q�1-Ǘ[�.M�i���Uw�)��W�}�3��r���#�a�羪�M�Y��g5&���SRi@����֖�1���]�_چp#h�������>R�D��70�t+�ֲ�@��JD�/��me+0���[�[��$���X��b4�I)%H;��D"n_�L�<l�KR�}V�.齼�����!fw��ﴜ0O[]Q]�C��y$�Gp� �SW��0��i��2h������_T8>	B���(tr��G��
t%��*q�9��qШ?vcyĈ���t��l�"Ҫ����{y��Y�[�kA�=��Bk�s1?�uo����W��K���'Н�<"�8�S�L�)�]���ʄ��#x�G�6��א�7o- ޢ_�B>`��y�/��~}�&����+�8�Z���DO�q�g��Js�$F��l�j�1̸Zf��QUyC�Ǵ'3 �a/�s�xw h�i�����N�N�&�\�pQ�,FAs��{�/�$q������8+�]TL���t��}�����D7���{�����S�&K$�h�a��+������4*<W�C��¸l�/�ZV�Pu~r�hr����X�+�q�{��n-�,�}c�:�FCMp{��3�_��%�������o�����q�
7[ݩ�H+An��e�JL���)E��[�R���ݕ|�r�5�}��3��J$Q�.�S֕/|�!c��/7J��E*�?@�C��44틊�/�^����}"����LiC��RLMu��n����SM���*`�YD�\��z���цy��W���#�eL�����i�7q�h���^փ��Ӆ�;����L�������7�w����7L@�5U5��`��ko���+��޷�7��wT4����E�3�NG�����p�}ͻbm+� p��V�g^v��*��\�]��|ca���Z�����#�B�Qږ3b�L�k�wV
COt|)9nE�Q�Z������3���Un�z�����m�3`����#���m�ظ�4Y/���d��Ź�'Iˆ�W�). L�]m�N��!����;��H�<�1���#��u����@\n��N�
~�{�A�g�9��g�U5�AF
N55��ӫ)�SBs�h�%��)a�b�R¨fҪMg
kO���M��&ˬ˲t���~�9���b�*�ǖV����������"�yR�f3%}���䲢����L��dd��WU'o�* �-�z;�����F���d�o���l�ǈ\ď�8�5����0'�����	_}����<�DA��Vɴ�t_Ӱ�u�tLp�ɨ�j�M��@J����I�X�D҇��Զٕ���?��F��1X]�֔�o���rQ:E���$�>Ү��wl��p�%����7�gȉ�&�B4�,S�;3O�b���I�/G#��[^��3s����_��X��.��ɞ���$��#��mv;�?|�+�(��N+MN�`jOW"���|�?�j�Tᑨ�ꊱr��D}]��F��.Y(�'fD�5Ew]�!�'_�g=�4XdX�������a�h(��1hP71
� ��_�}�^�H��qm��V�&W�p/�&���CA��G�������hn\��"]��>�0�I���#�o�Zި�جY�����U5��Q�6�G�a�i�.�H�0<p~u��M���jU4��c��｡���ܑ.k9�)�K�]�Z��ל�N�u�3��3|�ԫ
����P��_������%[�;eK�Ep;�kX���G��W19����\ar�+����J����>�h���i��R#`� -�x�N-�F��H��ϱJ\��������'V��}T@=H�S����k|���y��Z�-����"��R0��4��F��<[�wþ�]����ش��clf�`μ���9����c���iɄ��Jq�˽wk���F_"},#�zd��LZk�y�ئ��&�N��]�}wv��ɽ9�@����Yb=�"���:��h��6�W��}�I���0f|C7�>�v?� ���Lcpo�f��f�XAo�4�z�O�����Z�@=�{�Ga����<����i����L	鰈XP�l�W,�P��:L3DM�Ϊ�fC�TLÃ.�*����-������'h���m�a�s��*鲪b�O����ݻ�e�3����.b���.�>��'��.~��� ��`!2I,� ��U�6�[�` ������K.�	\j�׫�~aa`Մ����&T�����W��ຐ�b��c�6�h�Vr��>��]�K Z:X��E�{����մ���ce�����x�� @QB�Lѻ��ƾkP�`Q��Y`���Q�6��K����5l%ڐT�:Υ]R:�����Q �cH^�ق��Q^zƑ�̮�cD�w&�z��� �H��ڼ�chiL�qW!_	���yù����>*�%�P���5��H4J�&�z��r�8.�s��P��K"0H���v�UH�s�l<�![4��J��,%�D�m�{'n��&�Knu��H�	6m�s��lB=�T;�0<��.,�G�щ�zn��b��</L�{�c T�>���dk"6{���E*ȳ��&���d(�9F2�Ai���>l�� PF����fZ�V�s+U3eҳ��Z����`?K����3�,;��as����]���η����V���g�"��-.��l7�G$�^��1�z�Տ�y��_�G4���<F��`��»o���Vގ���?���:���mt���䤯�N�K�� �/�<���gp���Pr3>Q�^�Ǉ$~�JӖ~�]{��X�{UE�C�\9t Y� q<s[H���ENt�/�.,�mU�\�:'b�����D
.U?��w"�|��5��N�|xFw�uS��z�4�� ��$X��o��-kE��B7��Rߴ+T1��ԍv����	G����\I�"�@��yy�E�_��.t�U�X6{i��Y%������%�P��i�8��}��~�A����t�?T{G�����i>i;����%Mͽ�|
]f�*1��j�z�I�x�%K{d4�� �f3N3��Y�8���=���tr ��(6F⿍wo��T���`�D#��߶�# pfpJ�(}d)��kg/G\\��i�������|�
���T��G/Xf�4&�q�$���?����"�ݛ��z�������,z!�쮵
����"���&85��F�2����u�f�Naw�mb�+	�+"�؀�flڠ��A<�-sZ��r��,)|�&n�QD@����8�s!����{8%����*FC��u�i�d�&1r ���O9���9�[pP�y����AFźވbr�ӭ�i����EFOl�*_��<y���9N('0�j�i��-o��;c�觠�vfx-b-^� ��W9��Ö.A^��!b"�--�)v>��%-�%��x^%�Dt=p}��E�
w�Ŝr2�H��� ��ͫ��$j ŨΝ��ז��]YmA�3f]�43!�/YaJ;�"瘪�ґ�	�.�����Ⱥ��G9͞�<U�G�7(f�m�]b�S��Y���Ae�ܖ78�����߫��u|5��ڌ{H	�t6\q3��
���*bK>kc�D���6�It$�7�;ǯ��C�}��{5�>ID��?��פW��$��6��Z'�71CƑ�?��m�.e7#"؈�f�p=����7�rn�$:ՙC�l*�Ȧ�q
�;`9EA�'�&���p۫�O���V�{VY�G|�{���X 6vg���lQH����0*]�x��w�%*��@��]`�DJo\
��%���R7����1�S��A~���4p��>lA�|E��^$�a5�����j}6Y�Ğ�[B"84ԐfT[�FT��"��hҩ�����Z���T?�g�~�^Dl�6$E<�K�x1��]j�ɦʁ�e�-+��^,����G���H�ľ����q��h1�A��s�b���GJ>����Gͥfb�(Ÿ�xX擋��,��gO����@��ԍ����/VS�[�)�թ��m2c;�)8�qHe��������s�� ��Rm@*����vYj땯ָ�#�"S,:�pJ.:Jo�f�W]�-�����Hj���[��~���a�n���&��Ha|.4�c�lo}�o,���UA�ȴŨ'p{�:@�N}��K��4js>V7�2� �@Hmͥn�^&����傩˺R=� ��ˆ��n��E�ҙ�C��-=�{h�.\�t���$�Fp$���F������1�(���a�냄�z᩵i�^Jo@;9�M��?)��,Ud���($/�F]Xs���7���d�l$L
�'ksAc�Ua(H�w�H�JۮR	g8U����QpM%��Ã�U�B�*!���B/9��:,�":mҒ�k���q�Y����O�&mr�C����s�[oy��Q�����CT��M�Bރ�e���H�� b�9n��`V�ˀp�YT�y���nL]$�o=�y���9[����$�-i�
U�q���f�=��ސ"-|��^��H�{Ф���o�G:�uI�9���S��E'Z�zs䦦���^a.ԶAҌ�'Z�s�<�ҧڠ�y�(WA��zF0��p���m�v]Ԧ,/.�~�R�mn��褨�4�
�8��k�O\7��t��F3�!��/n��W�޹�J�O��/SE//��`�G������O:�����>��9���+�%�8�-*s�;�M%CӴ�65���X���
�H'����d���
�����q�Մ�������P2s���9{�}�s�]M�\�L{�AV���D��T��6(�š�<Rwc��ƣ�L>g���t%�\L�v��֐qs�>qrt2�s��|'�S����ڨƽ\���ymf}�>L��(-��nƂg���m� ����L ��O�A/�s̛��%����+?��:���5��û�I�H4L��e��t�о��{�7��_T��2s�ȴ�>ö��ډ��66^5���̭��n*; Bm�>���3�!�1I6z�����sh ��HL-R�ȇ����b,�o�ԛ@���QSn�۪x�7
l�P�+�<�1�<��f'�꺑�Z���
���]�w�Y�
	�X�`�2���3�a�q�3+k�Mb���$���vO"kj\�l�����<BQ42��~�h�i��-�-��`�/=0��y�y\~_���>2N^/L���G�mJSL%��g���VK�>1����H�0~�n�9���i���������g���p�ͳy����S��8�6��2���Lnc(MN�;+I��Ϡ��i�S�[����6��Ik�/4U�B�Y5��Y�`e�U��(6vv�p�1Neg 	���b�8YC�0�g>�?l�a��"��΁���"XI!۶�t4;�p�fXm.�`O�S�"4	��b��a�&4Y�u��Q��t�*���LF�Ei���#����r��R�mxny���&��e�Y�F�V��O�7�h�s`bQ>�����A������z���LǸ�p\6����+S�,.�VV���(��=�r��6��!{��6��'�>L���\�;���{=SX/)�������=X������I��w� �9�9詜����'�Z��'��ݑ��Dx-l�_q�K��mE��|�����WE���~%_Bk�R$aٯD�������fъ�`���l�x6�����&�Q _�,Q.�y7�m�����%��rIƒ�K@�\\�)LO���9{������U/�Q�m@����ך̪�n�K�9?�����QŻ����+�vm�
kԜO���\ �l��ֹ��d@�G�Y�]k��hc[�8��5�햕 �9��0�O�II�n� T�a"�´�lO����}V�Ss�')�Ӷ��Z��D�w���A���
�'��@s�d��+eK�ՍC<�����eG`N�[h1��Q�0a���sP-U�(�:k�)(�|�1W���d%$Vƪ�]ט�~R��HD��^}���0�~�Iy�[�8Ʌ#V=�
#e(�˥�?�C_P��W^�g��/�R5������ec�R�Z�I_��:F�,)�kb������A�L��h�Ң;�A��^�,C3�z����&=p�B4���|�]҃��ڝG��ߩ-��Rr��x�aGF�����R��5F��]ZщYt�.Z~���Ҍ��G0={��8�&��`�>�2���U�MI>�"�t�l�����E�X^:,+��}�z&�2.��̅�?ƾP�'�4����VP!h�2�z���Q�@�b]�Pq<�.�Rn�����h'�R����lݭ		�/�o�R�Q�L�����J&0�#NH�FA�~��<����5^��;�������x;�,�+	c����ř��?�*�oh'V�7T����R(\��ό��u��N����AL@�w��э�V�o;P�2B����J1_�
���и��Wg��f�����g^eiO�M/ND�}�����n��3~�G�=n8D�-V{�����@Yb'J�P�h��r#��;��lJ�A�F��qz*����΋��ӆ&/�,{����=��fJu���51�)�Õ�����!m�W�\��Xc��A�'?�'ä���޲�H��{)Lľ�n&�p�g�U���S
<��X�"�P���
��r�	�����ȋ��OI�H�)UQ������X��;�\�;v���� �'��',��Iȧ���=�����iG��H���vv��+]5��A=w1��,:Ѱ�.��!�"��va�E]0/�_�c����8������㰩��"�?�.c�<P�1�����e�mhdNh�qE�P�͓�t����d�Τ7�U-�KO�4��Ư�Y!����Jr�J�
�G;j��noq��𹫩_�N�i<����h^�=�����Ur+�I�X$7�:�.��~!j���29�Px]|�t�$j���!ӄ�Ɛ8\��)���S$�a�������JJl�V�MF$��](}�2ȮH	�(���҄C���:�"M���ּ���m������ft7J��M{Ʈ����7�4�j�?�(��Fs$�P�\���_V�No�g{r��	x/%�f���=X�>��}4��?~/����p�kˁ����W[�Ϩ��<�J�Zs�#��6���?:�jc���ay��!K�`!&v+�e�c�D�Q�a������!3�� �I���G^К0��a*Y<B2���22�����^�jeK����[K�*����{��vd��2C_��o瘝�So�=�%J�"U¥��m�c:��1��EZTp #L*(������.�(ʛ����б��[�Ƌ�ɦ�5mW�z&�_�>y,����cW �d m=;���LO��?��Ox��@�r%e�'���L�<�V�!ڿ�eW�z�#�y��b�As5�#�|:�,N��f��D<K�!�	vd1b_��X�3��|�(�i/���S/ ��@ҜFVJ��^��Z��O1�4��� ��I��e�6����ǳHr��Y�`k�~6z�JF˽�Um�O,8�a�9����-j^���!��˦�,��h,ook������*>l�@\�M��S�^�����G����U��(Q䠗��56�Q\4	{���w4�_[���x�x��X6K�m5p�)%J��nyw�H1+�
-��2 �/�/�)q zs��q�l���z��l�$>����V��~��"	#V�:���ο	d�9���X�3
.R�|ϸk��и�����z���ݹEO�e��#��4�ظ�v��M�O���A�unJht|�u��&�]���d�����y��W��'��/	sl��vtI�G@��$K
)�f�Z$�0���7;Zo��#d[kp��2�M9>}R�B�{F�/�Ƚ�Cb�'t�h��������\�BjN�9��<c�
�����-d���v6�Pt�8���y���>���PLL���D~�#��?�s�����~��˾(�F��S��[=���'\��x%��8 $���Z4���w�qu��>�|�k'"�u�Y�XJq�%�<� ���J��E=c$ �jE�X���T�R:X�4J���=QH]3o�Z_���ֺ���>Oǣ���cV�-_���xa&fJR�S-RD�Jr���-��e�c�{��2Ə����C��K;sC��x�o̡���'n|�"!(�D�N�8$���y, e��M_3��ՙ�A� _�KC�q�A2�5,�̶��]B��Xl�E���ţ��_�����t����v��ϣ���D�4*ȷ�:K�X������Nx����K��sI�<p:}�6��9�Uc�:KW1
������6�Mƙ�P�K��R��h��n��S��� Ű#� 3��Y� 9Hb�ᅭ��l�����@��M�����DX�D?��p+X��f�r�z����B�� Ru1U,���W�����:���K�|����uC�����03�m�-��~��^Ve�����''�؋�s;Y���o⢧P�5S�#���;߶YF�:f8\e��O�Q5�S	�@%�|O@ʻ���u�3�6(�=����L��,�s����(�rO�g�	��|(	�%��Ǟ�g�EzH�7���e-j���,Zd��>-K���6�jn6(L
}��:���u�@�~�A��)�%S�y��va}�b_�:���R�̝R��K�3��@�1���2ak�;�Y5�	hH9�߯I�k#+;��[P�;Qj&�>τ�4Q]`����.g�`"E[�|�N�n���WP�.�GeCmn���*�6Vd�mm�ւ.*q�vhS�Ӧ(��\n@�浢���q�i�iVe����2��>���h�bq�n�i%4x�br�Mdp��q�~�� ��t,��~tV��AZ�������-���7W�sm�g�F���A5ڞ5d V24 �%N���c�6�/r���:d���Z��R�؄u�ɹ8?6�J�?|�X��o�.�\zDy>O�4�j.F��DX��hF��U�b)}�W�w�W;�
R���U#ȳ�A����&�������()�~��vwh7-&\������QQ��"����4<;&�]8�F���e�����u���T80:]��<@s +ƴ�逮	} >B�d�U:�̿)%���RN��lw3L�Z��F��J����)d�4��{��(q��z��Qn�]�-��%a���/v�VHvJ���=:�B�G�{�
v�[�!6q[�u�Z#���.�?)o������+�Ӳ9�4�x�6�\�&N�G{����CV�1�� Du��P~�C���yS@k��;�m�r)�F�p�l��8�u�ކ�%���-���������ߗ�62�ѝ@���x���U����يu;s��38�?��X�r\�Am/r';	�n��;�j���x"��r;�_CI���Id@� d�D�Vt�0��~�v� �����PP�Mo��yjf�[��n*e,� �荠9�9�k��%����o i�A��j�B9_�3F ������z���k�m[�,�E�?���L��S��tv�L��%a��?)m�oe���2�Fl����2Ɲp����E�J�.��$$���!�.�5D�iw�˗66bK��ڍs�t�e1��R����U����#�Kf����>Hȼ~�_8n��+Y+!�}0&
j��;����m���T�x�a��
�WL�}���O�}I�,?��Z���"lS�Q_��I��3�"ěi�EM�G��g%�%�RA�[��?����ST���{�a�����;�]���1.��j���F�+|L���9X�&]#�u~�e���B�A �hB��s�L���1��Y��j��fN��n-��Y2T�Z�xT�"F�N�@��}���v2B��}-'|T��Ɨ[�����<��6'��t��(�{�+bSH�eŁ�23����V͍��>�M��A�����oQ�5���HLv7�_-6̞��O��E)�tG���g�kό�;e�J��&����/\P�I$=��%Ht�:�d*S� <b���Fin� ��Y/U��nQ�*��2 �.]��`���Ue��s1�o^-��t���]��p��T�&�vݫ��Xx
A����3���bR�1�:���(�0.<�+w�8i�?C�Y�G��!0�F_���9�g��QG���<T�LKI)*m�z�k���1S����G����{]'q�(�m�2�ޘ���JʘIZ�ʎ���z�n��k�R.�u^,h���r���p�
���BJ��2~�V>K��s+ţ%���Ә���Lk��{O#\�D��=�a�a#
{0�}zmEaB��sbsD��&��XoA��S�Ǌj��w� H�ާUk��|�R�NQ�Kf 30��6��'=~�q���iO�_bQ>H�$�r����˟v��r��F��OM\- �>(S�X��$0h!>��}D« R��(��/�oV��ؤ�e'�ʊ�p��Z
�[��(��=��_��2�!˘��I�(6.�㓔0��"��a�Bx'�χ�,��<���F4v�8P��G�pQ���1��#��T�/|���ER����鸘��\�|λ@�.wĎ��·ű�9�/7\?�_c�5}c��آ�\j[��Ӟy�	~��J�X!�j`clע��� ����m���eC��T��z�X@Ze�|����g��E�����x3��f�Y���p�w(�x�&�RQu%�$��%)�U,����*Ϻ4��)�K�,��֗Pc/W�6��V&+���j�e�Zm�A1ӑ�ΓN�c3��璒`J�x����h	cj��C �2_Q!�g��X�V+r�إ���jQ�k�R�#@��o����~��󵀅�?���<�k�dMW:��&
<��Ǎi�Bt>x���x������I��  V�Vߺ���1��6���Xn��5M�
DSW�(��c�Ej����,�C�������& :�&�x����=Z��.S��%K�K��[���\�ϳ{h��&�c�3c~X>6[��k{�I�$r}���Tȝi��-4#O��\����s>.$��T�g��*�qGO���'C�P�o�)��S��¼�H��n�=,ew�x�P���c��,A�=���S��N�^{H�t���4n'�#��ݐ�7T���O^�|p�#j�VZ��|��+�\R_v؆����rX�v�s-��¶Z �m!�Csƻ�)E��V�q����f��(���&Сj�����xX�v���7Q�0� 4Ys��.[� kr�rDG�R�P	RI*˯�Uћ����+D�%���a'�B��{s��_{y�]�����r�G`5.X=��T��6�\ˑ5H.�U�s���/,Σ�� �����#:#�ЄjҖ_�ec^�.u"q�;�8ȉ�Z x0 ����֕^�[�cT7pɯv)���ˌV��rPm���E@X���Y�.����X�I��[�厌���͖;��*WF���>�ͩj��W�ZY�P����D����hR�T�\����>07%���jG2T�ߥ7�i���,�$�4�`8,���9� '�ǣV[}Gn�3��;+eh������S��d���t���ρ����ԡ��?[��m�����C�lI����bL'qWO��w��b��8�(���u�`�@/�ݐ1�Պl��N�c~���0��R�&��I�D���]��|}8�&�QqB� =O@8�o�Z��F��������M,k�}I���vJd>�=Vd�<�I���F��pӴ�rs%p�)�&��6b��}�vS�E�o}�?���}s��ԣ����)��^�l���2+��;W���*��EEx��)"'��.���F��O����X(m\���7U9< ��x}�8��HL};�G��z�>��;>���9�#�U��I���@u��9}:=�	q¡{�Ϡ�ѿ[�ېh���)��<FA�'��c��=׎cH�ք�_\�Y�הG.l���}@�\��LȑOW�!�dz>C\@M���eޓGnV��> ~�JL����W�e�nO(�
�uǦ�� w��Gc�&���{M9W�"`<���.N���A�I_s���">!�ƴ���bm�q?����NU�����;#�ӡ�Ʀ�i���?�r�CD������Z�1��z�uy���W]�c����Z 3o�㖊U�$Ek�j�d7��i�����5�L#��]�\�Ԍ���Ʉ 4H�,����?Md��Q�t+����33�ٔw0aw��)3��5$=��sD�߬Sew�%Vv�`l�;����T�u�N������E0�u��ܬ��h��Fa������_.<���!V<1�D}��>0{~�U��q#/�Ӏc��EX,�b�M�ue�N��&��n"���E�<�t�d6�ᱷ,U�?ȴ�<���{��K|`�3�C��P��j)m��6{3]�����2#����w+�<4��qWG���"Z~8�7��!�Vcֳ�Z֯�m�$���;*�v2�f�� ����/ż�?���}�g\�f�)�@�FW@�*��1P�{7B��c�\;�C��f�f�-�K��#>hӑ,ݝBm�.���bngA�U��r��B����]Xw��#q�t�L�7�"R��`�t�7����
c6-y����!u;�f�ST�CP#�Z�\t��G/ Wfs*F3q�$ǧ��䖤u�$ ��,1Di8:<6R��5�U!ƾ/m�z�04h��).ܭ@�,�����|���噍`���Z8Tm�9��&����=
:�H�a;}�P�JQx�N���g���1�j�Y����4`��'����j٩��t�ݣD���4�?A�~���C�x��������1���x�X�]{����:���;|w�u�����wi�n瘧��X�9k���{v��=Ҿ��x%O~��u4@Q�x�;� ��}�x�$���^�xn5%�)qx�W_ZA����:���6�̄�_�U�V�{-�E�2��6	E�P��yT�o�*��)*��=S=���h�\�gQ����ڈj9إ�E��=['�Q�:�0�.'�l���z"y�g,Md�|�+���k$.#�)�Ɨ��zv��K]�]�4r��W������O�~B��2�S@W�F���ro������)eP���ZX�m�٫I�����(�
'5�7�.�5����J�\!���� W�|�o����|ҋ�-R�O��=�S�N)���q��}�I��p�G!�,���3�ߓ[��R]��b0Oz�������������M�FW�^b�t౻L�n,{��3�W���0F}3c��L���BpB��G��\��~�#k)a�3��s���9��N�`�-"JY)�W3�yx�,ȀĖ,P6
P7�#9�ɡ��ͥ&�>�"/���7������s=��?��'K�֒���?&0&R\�$�m��#�N���P�����^��/�e�X'���k�[.�e|�.�?�:_&��,.��#��K���c��R��4��x��l,jG|��<��捿��zd�TԢ�YL��h��x��`�+@�䎢��*n%kl���j �_�½,b���y^���+��@A{
iQRE��gp�u����{5�K-g<�h,:��g�a���Z���<�,9?|�j��\L;T5Yx��6���(d�
C=y��E�ժ]!��xo�>�c��X�ݤGu@��e'j�&ק�R��]u�`�	f��t�����{5o.���:L#�h�WY0}�폡��]��$U�pP�C*y��r7��i�+2������l��`HRX#[`�!ɑE�(b\p{�?I�52��U8vp��� �����M.*}I�0,�:S���}cU#�yG<&�&5T�V�\!�����i+ޡx`�L�,�6��O����`�y� ���5���Nm��N[Ҿo�R���D�	n~s�_ �fC��J���6�AG���a��1�X��[�j:�f" �ö������qhV)E���!ENl�jW`��S�Jȓ^m"8Љ+��m���W_��~)�
��F/��3s�(^Vh����ycx� "��,й����~�Y��i}uB 'ުn)��l�Z�z6�zl�a�]X$V���e���\�H����P2���e���U�������l�Q5�'�Ke��ϧ�ˈ"t��W�_!?F�~'V�^�Q6�F=��̷Ԣ���v�F�Qb�1^������z��̪�&,A�!m�{(Z�5�"^8?��/��x�+�"A�t5��� k�
Y�/Vb�Kd���|��nO�
=���G��)q��Em84
���^�cB�?���Q�3���&���H6-����ǒJQ ��ZH�O[�P}�b]�M���b6��w��Y[�J�.��Wj����Z�D�2ŷ'�pK��~p��HA}f�1�yu�9;�<��yP��蕣J��q<7�3Y5�Ma�z���0�(:$���V�p������"(��!�`����B#�,��K�3���l�F�0�d�z��)<����>p�V�@�u0	,�➂�Y��I{w�EªU�=�_#���^t���8FgU/ �+������[�Q�x�q����6�
�߫�v �hY��^ۼH��m��]F�g�礄��ܒ��02��p��Q�}߰��We�e{�^�����{ݯ�EQ�-$\p��&e?���t���Ak"�!�F�מ8<��v?Q~w�:��Ml������y��{���Z�A���s"��j��K���O�ԯևN�2�U��V��8���k5y�/m���5"ZYd��L��
N%f�.�ƛ���Z���;����	;00%Ы��٧4>�f�"�>7H!%�J�\����u`d��(�p�H]����oQ#���ꍭ�w��	D�<\(:��L&>�BOf T��"t_h��G�'H�Tn���1d��K|	[g���#{�=�pz)�\��5����RNDȜ-=�>Ӌ/�E���V#��V��"�r���x8������p�p��ʆ[�� ���KT�"�������w�V~Ɠ��F&}I�E9���	ui�l���q-"&�UN�)�_Vj���~{��P"�I��TLƀ^��D1��B����˛�N�������% $LF�c���	����*��U���f��U����B��nA`��Od�k��I��Z#�Y��uD"���g4��V�1p� �����ji��ښـ���Q�W�YV�r]G��DY���]��l�2��pzu��u�Xy�˥�:X=�b7�0�,���!tU-���[i�o�+���U�_�bF쌨u5��t�S��I��HH�3������Jћ�5��O�l6��'�P�4�a�ڂ�Sx�-E���>�\���[����%Q���4�c�1�>S��%1*�zh2���$9+S�$��F�v��R3i�X�����Ǆߢ��1�R��aӡr����I���F�I�k\.>�@�̀%{L.h���-0h}�e�%��uZ!�Ԫ]h�����f״�"LU����&X_i�ėZ�:�x�/eck�@�D̖��R�MY�͏����#�� ��~T�,Hra:CB�R�z��޳�#k�'=��8��f�/I�B�7��^���J �G�2���ЧȚ2=�d&��+����:�ђ�N�ؖ?��Ms<���El��8���-�Cy���6�xK�+���\}������N29�Wb��
H
��rj���gÙ��'�
UqK5��"3���&�~�#)�l����R�x�Q"��cm��0i�-�9U24��vc���b��TY�&�l ]�;0��t����v���e�Y��@�䆜F9N���l�_��h�E{���k�􂂿�:��]@�1 C �B�3��h�%��T�9Ǒ�[��R�;�v:f� $&����	���7��WwB:D��03���j:�$�:���}�xn*���J{9� �6�<]�cc�g��y=��X�{��U�.�t7k��,�M�_����c��?uN�/x1�]�q�YSF6J�)EQ���a&lCކf�K��B�����JP ֡��p��G��%�\�{���*���@��tH
ݮt
k�X��ZI������M(Q>h�����'������C�$�jW����I�� �Ca� ����ݑ�2�E�����T�-H���-��6/�d��������iV��sh�H���v�*���gw�;`�K���a�H���y@j^ϥF�\�찻�����j[A���9
�Lg�(VtB��y���kX����B"ث�3=�M��k�e\�k� �'�{.�;<\�WPr��FL鷺4�?@&��G�9)t�5��M���S���5i�1���n/�\2c�~�Lqg�*`��'&���Ӥi��mMv��)O?(ʥ�F<�V�.�!:RkIa��BR�|i���N���͞�Ѓ4=���tÐc8��97Jq�=�����o�}@<՛�KC�}$>��e��s�P;���IE��=�i��1��rU��`c]��o��)��#�qw�#�~�~�ql�C��^��l��N��7����ҟ�0�O�X��<�-�#S�bW;uX;)�)�a�\���O��� ���'�ࡒ7����M�������d]a|�lտeߊ�#�Q"�|+49��(N����m_=W���{l���:��������WǱ�(B�S�L�>U���Z;X�ЗM?���IU�H��m� )��0`�O|�4�Qs�c>�^Y��}�� c����h񯉲RN�K)��>s�[q_)��������؀��`M8D
 �<�e��h�A5�A��s�M��tΥ�T����{F"6�Z��,&ӷYJJ8�(Y�!I���|�YI����1�����L��hz&����J��x�>R(��#`v��U�)�"����\oԫt6#��+J�t����?7'ȫ؟�du�ե��P��s�2c�>0"�sp�A��]m�0�ō$Kx�׃56Bx4�6
<_�k��0���ο��ؕ�x��d r�3�B �l}�FP�"��P�7
����uB\ ή?N��a(����
���S�7�Hl��n�L�)���u��~��?����B��F�+g?WX���� ��w7q���1ظ�Vd�T��F~B����z*�U.Gh��\>�*^�Ya���๹E!��Jm����U�� �Q߆�L2���f�{�Zb�C��eR�1�������JY�Q�?.�S�-��Q��T_�:���'�@���1����̺U��t�ܫ�$�N<�&��SCC���H	���b�4��(�<{aյ=��r��`�DL`��2w�G
��W��O����M�r+�>K��7� cF�����R4�>
y�(iiI�`T�	�W��`�
E�)�l�x8e����1��7��1�=�:7�rNEE���u_:Ln�l��\#�u�� �����'Sw���RǴ%�~z�M��A���߯'�e��lQc@g)��N�*6���ӀZ�&�m-	+���m���E0���@���f�ʄ�͌�i�
6O�:����hgNQ;(��������c�i�n����x?�l��A(ݥø�~g�l���;��A�`F�2IY����8��q6i#�u6"�"}g����;�������qtqo[�u�ѫ� ��SB��VݨY/}{+��wJ���v(b�`�KW"�_��<�D����&�+���+о>���6��e�T*���RRE��U(iOi����qH� 3�g���J�)L��o�[�X�+eȡL��.3t
�c�l~jd�2����Ԯ�Q��&�-/k���M����e:�GC5�X��i�J�~���C;�=Zh�24\�m�(����<���
�����p�x0��4 �;� or_�0n�]f����������>�����.��������j������ѿֳ�e8U,Ŝ�`	�n���o���/NL8A����;ڱr�Z01q ��L_ �r�����$���>q��F���j>!�e�ݺ1b���p�i]��m�_Q?�dR���ē	&��]v3��-�{�5�e{���7�g��Jv�:]y&��<��3N���R�06����@Sې�`�Q̩,�!���ȭsk5��]I�H%J��;�F��z{��ev��@J$��L��1������Q԰ƌEk����cY>��!*�o��%���������	kÉ���N�29� ���������i~`����&�1�h>1 )v�D{�=��/mˍ�F¹&mP�BFIh��ųt~�3 �&�n.2\�?���	�9L~.Њ$f��?��%���Eۀ��e�F��4Eh7M�v��ŉ������7�B+�w�"#����g[��f�#AFqR������r�y��腺?��*g��ѽ�q�~��`�O�l�6yG�>w.�ӕ�U6|s���l=BLQ�̛8�0:�z���{��#�T�c���eLCN�d5&�MfcWOq�:�ݤ�����uė[���o���v���jSL>�w݇M��z��d�^�u��!MU���5=&eȄ�d6@������!�ʷ��Ww̓�%f�E�	�R�:��U9��������x��G����ꁷhj)>0�'�Cg��^!1K��O��`�[����^P{��Vg� /��5��Ѝ����zm��hW�R�|ށ�)�ܪ"Mx�<Ҩ?ۤK6q1H->� $��Y���7��ݴ�v�t�Bl��ڋ3u�19jI�����X��@]e�s(ҖD���L�u���	}7�=n1M�V�s��$�ó$;��_	z�(�Т�-�-�+�X^��!���q r�>�	3k�ʐښ���t�V_�#U^��dCd��1�ש���Uu�M��sC@
�͎-e+�S�/k�!}�~��#�h��[�*U���1��ګq[�0H��}9�&���z�
����n����U*��bY���.q�^;`�/�f��mf&�>,����g��-F<g�=�q/N���t��������Ş�<"
���nM�#Tz6�?[j^sd�]Z���L��q�����U)Iw&�g�hG�'�$�B�3�~��&k��H��������c���Aw3�g��~����Z��ϒ�K�1,�;�tKhj\L����,�}�mm���/��_g��(:?�G�����s�S���s%�Nظ��3�g�����뫵8��ؐ��#@�����Jd74"�Һjr�+�m��Oպ�^��M��Ȥ�w�����_����J���Չag��6��'��%�J�n�0�
����⃰l>o~��_��o�����W�x��S�x��A3���珡ɳ���A�I
�o��Z_����ё��';���R�B<�De�� r(��ݜ�o�XA��}��� 茄y�)!��Ts+�D�W�����Uh�8�%�4E)��<�!O��h����t����]�x��Q�M�������!���\�R`c7���{)g���M�� J��w�p�A��������60W"8�a���sU�9�,ت��2Q
p����0H��@���A& � �ϔ�՟����ܠ#�#Y!Ό{��ˌ���	Χ�$ޒ���Ba�P��F��zP�,�x�M�H�۽bʘ0UOk�y���ڪ2� kWt�A@d;įc7�L���D�N5���֢p�-�3m�QEPr7��_�X��]uЕL�B�R�w&9ň���F�KB2�Q���
m_3aF�&z���֕��dB8$��H��-�`�	�,��phvŕ EE2:g�T��rA%g7��,2��)�CN�d�N��Np�.p��'���44�����Hi}�	���&{�rC?��`b��ĂK��KV�p��Š��Jf�3ߗ	]Tl���K��%*f ��0M�j�[?:B�/��SQ��x8��Ŧ���-��n5��X��"'�`����ݷ@N��{P���Z��#nR��ҝxh�_cS����z<Y���bl`�c���>��Y�����&���:�X�[.�D����C���h��y���s�I�ADÅ�_�5P	�
>�}X�eg���Ȉ~kM!X%ٻ���c΀��x�U'c��ѩ��U�*�1s�E�$�trd���:Z�f~�q8mt���l�,���x��pb����&J�ޔ��33�������n�HU���K� >SpR3���E%	V��-�
V�%��%%�e���P����h�����c������9���u��4|R~{@����ͽ��U	}�:W�vp���^��2�]	]i��dr����m��R5������[\�1��!�Sw�ӽ�a����������˴O�S2aV]�1S��e��;O��?���>��5щ�TN)�$b�����VŴb���6#��˃�4D@(��D�=X�u�{{A{�A��|���)�֣i�p�A_@IWa��hgV9^8��?��8�$�m���Zs+��dq�x|hg�0ϡ�z�>zY{L ��1�x�3�v�[�Q������'3\���+��Z���+�c=�M>�)��Hb6�=��D���?����j�}�&_��9���U�4~bvj����9�0�x��ң���������^��`���s-�3����`�����Fk/~^��N��qt���ur��5��J+ �aB�R[�0�\C�3�A� �D�pS�'�W�޼��x��1���/����
[���Q�C�|�a���b��AzK(-8��n��N�.@�'� �D�}('�3�j�PIBӉL�q�3;_c�O�ܯ��}�"`�.A�&qn�ED�xx<쐪j �]fBT�/�z\�M͋0On5����̵%�+�Ja�,lX�� �W,��I���>�nX�%jD�q���[H}�GUn�cR����fR�N�����Ό���]��O�؆��@p�S����9�#��W�S	>��sQ���Z��.���[�c���w������|o¥�_�4`��tԌ\(Ը��Gҙ�S	66�H�n�r���9ⱅ���|<�ʚ�\�u�6o�=P,�7������W��I���Π*!JZ;m��S�E�Md;�5�MjS� �����3)�RA�ru~&�H��-	��^���'�����|v��kD0���'��p��J4ڥa��b�
ʗQ:꿉��:�3`��ظ,0z�#��	��%f��[�5s�Ϲ���X~*}LB#�{�Y8.g�H�����I������1�Ě���)|TlӢ(��&ʇm&�R���#�c�)��8SLEֈ�X�T���y!���a�9wc�wh�Ѐ3�����|ŁPa��-_�;�G��pF�i�,{�K�J�ee���r�|e���	��Z�nh:�<&_�+."'/۾����鏿J����~2A�=�dA�yt�̤��QSl�����Z9�%-�Y�����DQn B]�/�:v�����;��O2#BY���\g�^�9��2����ս�tX�OH�d�s]�d+�HV�%�x�(��1��m��U�<��uЃ
�6�ҹZ4(���zw4����u�M��j�6N�*p>s���z���v�ܖBe�)�3N��e��z�""�T)���rw���|��\�_ӿ��w��S2��O��O��)�ieـ���
�h\��7(~���@*� ��`�EbB�0R��8��'�Ύ���#���7AH���*�,5�sLΣͲ��1�^ V`�FRw=�B����r"�?1ب��z[�a�]f�Z�m׉4�̤	�`s�5�{$�~<A�)'�#�A���{=s�Ӂ���?i
�����J�IB�U��nz�3e�[�ܛ�Hj]Y(ֲ�,�ܺ�N��M���o0xW�>_X�W���i�낑��#�l9`�X�m�<��㻞��}fS,��坎e�L���te�IY��O��2H�����כVz�l`-����r�\]�v��r )9�hpB��[�N���bӋ��>�ĉ!�׏�*�3[��;֭iJq��21���D�|5m�q�\ų�F�X]�s������1�n&J
}&@�F׸7���Gg?L�.�p6�s8H�/���V#�SUKʑ�J�Ƀ��A6�����'��m�V�~�:�%�I����yA���9T\����H�x�b�2$��2R�E�.!�%F������/��C=�sqW�FMDՒc<����]�y_�$�FeD�ζȔ����
�������\���������1,�'�&�"4
:3����FYt���:�kmNg!G0�O���A���RE����B���I��W%��d�����a��Dg������יNK�¹�]^��$cg���Y������8=IF���y�禗�H�%5�O^���)N*(�8yI���Im◓=�d*,\��ü�m!��)���K����)'�vGL�-L�,���" Wyﳧ<��0�=�"F;� �����y�EruV�c�����I�|L8t�v�ft����!�i��/}�����X������V�@Xs/>ABͲ�0��0zMr3~��u�~����<G��L�,�����ɾ��`�RC�JM����8�x��`��нV��ݒn*�v)# ��x�2I]w�2<TO�"4ZJ�BG���)��7�j�{R���Y�j�_�1�����~d�Y��C��{�Qd{P�8D#�f陴D�5���#f��'6o°�5T�䶃���6�g�2����q�
���T�
�6��S4���cgi�-��\�ٺ�K�A��cˀv���!)nK�2��X}����{h\�m�|�6�l��W3��#�3!�<����خFQn�t��R��$���EU��V���p�|>�Ӕ���R~�����J|n����؉7�;���E�~@ҿ��*�y�,�ť���t��2j>�����m{~�X����Oc���Ł�H��$�D_�D�(�g�Te��T(�]�nR�t�¿5��&�b�S�K�V�}���3�I(�}���G53*RT���DN�A�7˕'��^���@������ H#���@������4��9�_�CC ��p,+/M��t(jA�(�l'_¸a78 ��9hN�b�Ѹ#����_��3�K��c�����ו�B{'"��z�Պ���o_M��-ds��e�������P���(+�Ԓ�02�^{����h��o�Q2Y��K͂�B�SAQ��/�QCҽ
��Y�2\}EĽr�>JK��j���i��a�v٫��0T�	�Jz�w�A��q{���<I#��8 �)N	�� ����Jb%|}�|�r���d_'�YP�/X�0�Ϭ���N��������t�a���L�2*C����ײZG���%����ӎ�R|ٙ���g[TxH���	����J�D�}�ƔE�G�u��+^�}H�_ҷVr���oWQ2�
�e�.ҳa;�P�CA�!9#"&(���`S!��GH3�]�9�̗֫�&;������Ź�7��H�	a��#g�Z#Dx_F����>�+��"�VH-���p�����d�x��l3��ڢ�hQ�Ϟ�$��(�
�q�k���C�G��#��boN�m�#K8!�=����+�bRcOH:l�Ш.¿�9�]������� �m��9��v�iTf��ɜ�����v���p��iZ�`��S�S���Ь	9���B��l�7����A���.�x�U�d➹����J�rf���걛��[�O�TgTy�2_y�*� KO0A�3eLi} �헆v |J7�8�tEj���dh���1~B�p�&
����)�h�wm#�Ē%���{T|a��C�G-��W"�	~�yql��e��JEI��n�9K����ml5�g4r%�%߷�&8����P�Z�4���ѱ��HC�bg����ܲ=���j�14�}|qz5qd�����_Я�7�\6��'y@���@(����+��b��C��	�t�!��d��Ͽ�Ev��]�g�S�n|%x�����9 ���풔R��_��|U�O{��@_ཤ![���G ���]DQ^�ҍ��ha���Z�[�D�����+���t��˝��tdE@�kV#{ �e���~��T���O�	܋��p�	�'R]Չk�No��'aR�}`Ɛ��qV:ԲD"���_�b�V�0�n|G��#e}̀�fE��xUǔ��/W�4���6�iD��p�]}�4��z�����8p�Qv0�,=㻫߇qY����*IX�I�є��_d��Z�byc�C��}|Hf0�ȇ"�0q�~R��PV���S�7Qe.����d����;q�)pj������h�f@	4��E)�h?7�w�)Y!?��G.-���.�a��L�ԯ����o�]�q�Q�d��Y+}���mG�uU���{r�C�(�.��p Չ�dk��M�"���?)h�>��d1M��ER���o�Т��p����b"�Q�C��d4�sO-�x*�zC� }c(X"�)u4ǘ	���Y!�oN�uk�4Td���KG��4�t�����#Bgƍ�d�S�.揕�;�{�$n���Dٵ��Ὠ�yHyT-ۮ�O�T����!�U����	��0�.F�
~���=��Y.3_�� ���|m«\K~i���P6+�L��h^O���1���[�Z��fYB*�B�sy#I.�L�(H���e80"�H����3���K����`i1�"W�'C�o�P�U�}��w�D}վ��1�}�&3�-G�3�5+�,=E|��d��)r��:}W%
��I�έȱz��Y���t}��Pk�;���7��"f��+�������W�i��tdK��-Uyo�a�:����
3f��rg��H���ҤR�@_8o�1��7�����oc��v�����S9���w�R�ꖭ� ��$4Y5Bg��q��2C��%J�Li�������"����W��2њ�?���ц����
�����Ǩ���{>VJ�<��Q�yu���f�Z.4�el�,я������`�M�^��}�=[d�`�y�[�J��%���u��tp��\q���L7 ]Xɸ>A�$��8�����h�3�ҹ0�=���)3�!M�T�>n��0�9�������¾�j���2������1#1�`���Z�q�ݮ�h�"K`ջ��(�y��(ÛlU� �6m���KI��V��*�:#�J����; W���T��b�ɘ�h��0�P8��p)�;)�o��M�v�'�,�1��H�"�J^�'#�H1׮�y�y��ŗr�n.[[�XYa<e��c�XxyZ�2�p�ai�>�('
��ļg��r�.�ʰ��w+���t�ݦn����:(:�n���Xj5}��<LpȪ{V�C��LgG�� �R��j������d?���ؕ�`M���9�ȣxQ��ǹh�}��;};�4��`�t�q�VblS,�sQ�H�������(���'y�ޑ�F�	j[�
�5l4���5zH��>.E\%�U~ӳ ����T����_Px S0+�Ja�>��qb�����-�x>�'�P������]�|��gw�˺Aнq�$V���?�$��׳���Fٵ���S���p�[���MG^6��n�����s�	޼��=�FT�� �$�ʅ��������VAS��I�ϵ��Z�xre�P4Y<a�4���=1&(�T9�.�g��<}qvH�[���ֿ6����s.��Ǯ���=�(3']�&�����Ey�_��D��k4���6��m�O1�r�&�����[4�?q�(��	��lt�F���"�9&s� �n�Ls�Eu#TR��u��MI����U���:�DrLNe��2sUh��~g��.�����m
u�o�q'��ؚ�,���6�����XV�dX�e�L�\ɕ�#�Mcl���w\��z7K�$/C���2i�'�uN���-ZI�B�hA'��!��q�#'&S��v��s��H��z1>�iI.TVB�~D-�?XW�[IOH���νX��
�����i6�{���ſ	��9ww�� jq�UK�n���2��d�����Ka��tv��-�y�0�2���I���gLh��5D�t@ S�3���~�ǃ��K���}��
;h}�E��bh�T��׶�E�K��Ӟ���8��o��^p���, k�4��Q1_�J
�ρ�V͚��Dn�"x�ƻ�_b1o��7ҵ�D���7�@"�5�H|�,�|ٿw3����G�w��-�P���q�!�|+��>eEk�oh:'	jQt��=gͣ�DQr_�Uۄ�k�\u^��4���j8���Mˠ1���v;�B�ZL��Q���tn�U�r8�����F��<���0]����M����Wr�O�ゖj�\5�(�8��%S'(�'��!
����ph^ti��w+zE�c�U�tߨI��$��S�~*KYU)7"�O�#N2���4%*y�����~�ڕ�ێ�[k8��<F4"�)4�h.
	�?i��9;Q����2j�;�?XVTj��rdד"2�WC&8<vi1��L���H�[�z_���L�+jb�x���2I �О2P���3J�=�x�_4��A�5�}��6L�F�|���`M�y�ܵ��[�9�̀Y���3z������N���h떄�,!m���S2m�L,*���v��k�9A.��+�c�=�_������x�tg̜��e+�����Y/,��/��z���I�E�3��]>��7�I��`���~r�N�/ޤ
Vڼ�X ���/���Gw���R(K��@P��mP��ɻ0��(�I�A�(>,q8�S#G$�� �f�Xp��������Gb����K0�&�����GhM�:<;�6�@r��K�\#�y�&���N���� ��!}PFh���IHlQo�q��:�c4'mӤ�	����''���~���ku���RG��5(s�+���#&��C�F���0R�w���E�$χl/�H�a�=b�� 6�3l��j4&H��*k�^O�D�H��Ĥl���~�k�\6¡T@{��(j�D_� �����d��nA��Œ�3�"ܽ��0ɗ�o�kz����Ƴ�w4"C�¸�D�����1�&��6�VM��H����~e��<Sp� XAیe�~u���J;39Zy�6ߐ4 ���Gv)�z(�H�$���K�_���_ǩ��w��1o��+E�#D|���W��9}G�闕t�7r�{;����\�Q��s#�����:��N�7+~1���P�{���9L�0�y�Z�RC̥����_�	09�\�[���!�����l5*F�l��G��k���FB-4��v�!3ȴ��\��|�kXYS݂4��T���Jv_�Z�����Vq�������˸��'�
��Cv$�Sөe�g5H���A�&;��1o���&\���e\:��^�^�1�!t�u��Rt.�+��a�BY��B&֫=���Z/&m(�Ĩnw�|F����u����X�ePe0�F���m����P\4{B�n����}-���($S-i�Zp������ �?_�g�S\t��l\�����n�H=�ı��|J��d��@fғ���}�З8�������#�'���(�DƒÛ�v����$�&����+�>>*�Ɉ�ܑMF��)��+҂ţ�W�$����R5;E���H�<����"����*��ea!iC�J�l����n}�r�]�e3'���Mh\��q���*��1)�d~��r�U���ER@��O˰��2�o�.��xJ���0�����i$4�;2 <���M�i�!�-+F��oe���;}5���#@u��e G��qd��3M~��u�2J��~�N�	N1�b��ê�լ���:׋�)�X���?��j�&�_��MY�x�_��q���A�X��Qi��qX8$X��5�$�/��<��`KgD~�ns�O��F%�[�y-D-L���(�Uܖܔ)�T��^p�]� ��H#�Ta��4��&����Drۣ�SE��A>GΦJ �YVξ6|�J��b��oWj���*U�����j���)�����SsQfci|m�w�y?G	/�w1�s�f< SӍ�^�Ǖ��99��"��,���G���4�������T���!֐��[��o�!���L;�]r�3ߓQ��d�~Nq����L���'q��_��w0+-�z�����E�dT� v��qU��˼M��*ὑ�u��9H&8��$�Qۣ1_��A!��,��H+��,�ѕ�����OLo����oe��d\��~�1��s�I���mH�q��gX^�E[e�#c�J �o<�m'�>����ش0�iӲh
;�����CS�rP�?֯�6���=%�nlx]�Ym� ��Α:�����!P�t�L�^�~�ou�NG��إ�����mr��U<%5��}=ڬ���D��k�~;0�>���B$����i$�^�b�/���LxX��yP�7{8�z�&{������j=5��Jq�@M0��R6vwQ��7�=.�'A��_44���cvpp��]lMR�1ěmj�b �Z�X/KBYP�*��A����<�N���U/���f�2'���<܄��o�c�T�i�����fc=;}4V3Y�J/4��@����H2�r颽��A�Ѽ��sa�B��^��ِ?�߷�l�=Ao�,��0E�rm�9DO�9Ȩ ��8�e��ؑ�8őh��r�Q�("�w`�����^IN}��Z�^R&FJ�Qc&�76M��`�v�ضY�tP4�w#L )��oW-�q/��9�8���խ5�"@��=/U˻�E����2P�ӒVZ�U����7�f޿9I|�S��	5X���k� 5_�q;�/6����hw��Q��s$6�=5��z�>{h��Q�J���_�f�Z �)=I�I��5	�ͭ}��M �Ά��`O.7n]��	ᰬ�������]Yq�R��r��c�\��,	n�m��I��*��88&�Sֲ�~2A���o;��m1Mء$[���<6wQϊ�n_B;+��;��c�T�{�=�7S���h����
#9Z�����VnOTZ����?��&�����|������E��seV��ν�΀1l�"��to����Q�3����Y��^��ױxT��D�$�e1qeǰ��� �խ_~�(���ɸ��|��r�}Dv_�S�F^dWKD��U�ȟ�n��	&�l����<�rbAYf�oD1�'�Wi2V|�d}����q��,�r�>[S�E&,������տx�mP�1)��5i�x���>2��`��٘+�rX��́D46�L��!����"��dz/������	Uǃ��}�0fc|��"�4WP���>dZ¥���G���z@2�dk�,����%\�K�|'�Տ��_=���'�ڪ���d��2��|�#G���b�X(��k�ݯ��`G�9Rצ�W������9v���K$(aԅ�f�ƌx�Xd��6���׹Hx�����Q��A8oKz�e66!�gׂb��I�����;�����(ob���K�]\|p�M��4���V��:��~,|Ou����
k��/�o +��I��3�0��}$��2�A;u�n�G��|
��4I���ħ�pk�9g�}Z��e݅*�5h�}�j>��ٸCO��mD)�L�����8��W�]�-��~�!4���s��Y�����>�k������b[Տ����՞){C�Z6kr���B-ZX��܈���H����
�O�'\�HYy��a ��ѹ���h<��w�l�D�(��M�H*~إ�a:ۍ2)"�$qhݍT��}m>�%a���_|uU��k/��a�&_���%��O=�"�x�R+ʲ��U'��.+�,}u�����&i-�7m��gU(�WC���� A�+Q�Ky�6k�;��%�O�S9[�;�	d^M�_��I|��I5��`̛��1���_�,K�>�7���2v��+�*����]K&�2�"���Hn��$��fA��L�k>|�s��<G}�rd���QYuS�P�h��L5�FpN�����v(��\�V���7E���s�^��Q��p�P5���:]��'�i�2��
X�@.4uđ��bѥ���e�~���a�Շ+�l�ec�lO�A��#��/ ��mR0��SOz�#�2/�~�?;&V�gD������c�[�HK~����ϛ�XhO?c������k���\���a�rc�ok�b���r�2+�Qʥ���b(9�5���,�-KE��T���d<��/�%�Ə=pj�2[4�=0���E�f�����=��;Ì�0���,����U��c��W����=t����fS�����s�$1�-�Hޞ�b�4���&W,���LQ�bʶR�l!�}'^h'C�Y$�����<���+^R1��ֈ��5��ٰڶ�-����C��A(��?��LR?�\gW�����ocgD�x
����q���0:2Uk���6P3�¹�Raq(�,�����ȿɓ'w�����Uo�6ӛX���(^ޒ���t�	��QRE^A��,_6��F��ְ��V\	�qk^qf��HA+<��i�T�� :1�ޤ�<zT��	�-�_1l� Zj��H��6�7)h���I��J*��h�v� Ò��Hw��Ib$Qt~������So�5��oB�`5ҰS�4��8faz�z�_]��������x!U29��\n�̶f��o��}�V�Z�'�I-�����l~Mz�lVj�;��[dd�щ;W������b�)�
�@]sn�0�
�_�q��}�r��M����2�r�C����f^�a�N�rV���t��$ep�lq�b$-�����[�,]��T�G�Ͱ�X=�=9�tx*�N�7ތ��}�ri �m������(��$Hj~*M��<���v lǲzewwJ�����Q�g�S�F�O��+��U��Y��(����T�\ܕ�h1��J��Ĝ>���W��I�%���C�ū�+ٕ+��(�����T�\/��#E����>X��������)�u�3z=S���7ϺW�WO�[Y��ʉDR��F��p�ز�o�Df�2��%����И�����0����aij؉��;�ԴLf�w���i2�����c��JG��)�������ꡇM���\�W�.�
8b#s��
�sa��!`��M�Tp�@ԜJ2��J�f�,SF��Y.<H�m[!�ג���#�� 2ҋ'����vR��$W�^F�O��TП�0��(�%!8.&�-}�1����xV%�
δ�l����TP�U�$����D
1|�����Q�a�����Ks�O�,gf���;
$�E"_���I���I�������ߛ~��'ߩ����f`-]��ӹ]��yOA�1u�4l�$_���Z?BRZ����'쮂�3��
��v�'P�cՂ�W 
��L=�?j;{��V��O�X+Q�t�A��_IreO\�3��D���8y�L�V��;��(c�B7�w�Ad�ݼ�@������m������C�.Ϝ��'Q��D�T�O����}Af�c�p��b6�|�b�}�'�Z�H�����5��T�S���#�ce�R��=y/}���M��o"�f4&	5K�u4ڈ=�F�k�$�v�"���qg�B��s�7!g-��Ng<ӓ�\Q:޻��hd;Y)i���j�*�`�kF�|o!�A��t#f�"<5>~�t�ҩ'�6��x� c'�����\¥ 7��t�珉LM}�|V,�LjH���0@�OXe��x�43�$G$TCq쬎���|�g��N�`$n��`�ESѹgs�K�|9�!�]i��z��^u�~B�~�� c`NZ'FH�G�A�=#ٴ԰D����n�8xp�;$���X�B΢#��Q�C3����P]���4�� ��O�3j2d��G7�d{eGƴ��ãx���e��xg_G$M�u��E��z���gxV�2��`+p��+p�t��tI/���ٹ4� �g0�V��}��;j���m�&�fk�ԓzB5ꜿF��m�~�NOGi�J<Ʌ�.	��0�uX`縲-ta-�?����<	���k!�i�ߟ���/4�]�&�,��RfO��_�-�R4�@W��TB2�`ԇC���N�z|��P!�/8$4�-���^`���.�:��W!�b��F3��®�x1@�A�W���;���G��ˇ�oe��u
t�N[���[1��*�0O0��.�K�3	*$�z�w��%/���*)�����=��g�e�Ph�!��܍�C^�����cǃWK��*���`Pp���:9~��z2���;��j�:���W���-Z�͒)C=��2����k����iPH��d�e ���"9*�k+H��u����h$u�m�"z�$%���s�n�]K8�D/E�:M�ɣ�`H��3���D� ��ߦ����S]q`Nν˅iD���]j��|ΟiW^rķjSW��0��b����]�eCx��0�2H-X�}?�:�C���%��a.ނ8N�~�[�]Ɍ1���U	����}�	,i0�,��Q�����[f#�Pi��fW�@Vh��*��/�7"��F�-�s��﹗3�3��񄷦A����[gQR�-���Xj�=�3*���nq�T���̫��/N���&?w�1,�ch�\Y�W�Jv�	+|�Y�}��C]��F�ջ@�C�c1�\n�j�a{�t��t��G�� w��0n�����13�&9q��FX����i26B�PMk-�6 z�Y��o�
gԋ9+Ou��՗���o0�L�EX�TC�j�~�$Mb�fߍ�H����G݂�E��KPE�5�����pt���0᠘�5��� E��,��U��O������
�>.�i'�L���5p��2��29�qz�l��d���p��Ŕ�E܀���]�����u�-��"�Ѡ�����c?��U�s�:�;�T���<:y�8�'j������h��n�0��LZ9�B�/��A̧�8S�y�q�]��<��e���*�Z� ͮB2���õ�QQ��al�.�^g~ܶ��¤di�е�� �=��E$�~~P��s�9$�K�0w�/�1�n�ڬ'2�Ֆ_�M�8!��ULf�6�Ng餂ـ��V�:m��� 5`lx[�D��O�W��.�*�ȃ�\Dn�(���ǀ�}��.�5�Q8, 8�WIаb�km����L��PW�:�(+.���-������Gw+��N��\�a�W���l�**�2���������}��e�	+^���/E�T}I��O~����6�\�2܀D�ؓ/<��I��G=X�b���]�F�~�Qn9�Yzqc�:Q@u�SO��i�	g �7�%�,�SS��u74�srN���� ��H��.&ے�ݏҿ��y�>iX�0�	� &pD������ʏ^��[�G)���Y�y�'�x��<<�*<���RT�/�~}�j}�	���D�I�4ᐥb6͋�#; ۵��H�N�����Q$���F�e-�x�V}E�z���uqeQ7�1����V��O�}��j�o!�x}d��(g�#�Hs{���q
<k���w�!H�ݴ�F��gp�|�UNH����h��O]��d�N��]��D:����j�+����Lyb$��S��Ģn����@Mg ����x�ds�+\�s �s:
��t�~�Px�='ʡ+M}��i�w�;2���y�Q�����g��V�G��$ˬ�\�=�(�m��i!�s0�xL���xV�(֎GH�!s�}�5�r����a􏋿�r��U8��kԓ��'qKҐ�x�<>yL�D��^>�]r�_P�s����i��u�mi|%(��8+�iy$����ry��c!I.���	˹�Ɉ����A`,:#�&0��Q�U��Fg�R�6���P�
��&��������-M�M��֞�
zc�K�?�������_�_�|��_�ɾ�p�I 8T��ETvќ2`�I����-�M���~�jt�O�u�k�3�>��Wa�����Z��N�2�����OȽn.�֝�W���5�~�a�g;�kk(�$܇/��nbk]�D�]��um�S��`��(W$�����eP������p�$���$�b�r�a,�7��T.��`� 3��n[��p�	�Bj���k��w�館&�����N�R^�H:�cc{�H�~�":��a:JbP��Lz�1|���Hj8���ɮ�p�F��Mw��[�-�҉sSm���i��D�q2�V��O��,h��车�^���K�H#�&!4�L�* ���0�� (P���~Dm�FD��W�tmҩ��x���k�'O����t�,޵��'o
�j;!Z��t�/��� ���K��o���z�gV�iρ&qƞ�ˏV��5��E�*>0��W?��3z���M�'a"}���hw1��V!e�Y�oM���P�Ir�[���7�#6��_�3�j(l�E���S5���\E�?J�4�܋��zFU=N����w���}�U$�5��z�)\�a�K��FTV���� �h}�L���_��/�U}����J�c����v�@�v�Z�;	#jۏK ��d`�5'�� �Z�Z`<S]*Q�D2��d�����-�`�m�����:6��M�qV�q��ɻ��_�ޚ)T_)�#��ܕ&��t��r���)r���S�_<�7L�%f����?;*Z��m�m�r���ҙ*��dm��
����lE�"O�%G��/�)�� #�lV�Yz%�W�>Gi�1\Ŏ��4����sO�R�=R���77�d`e��|����\Qj8G��%O��|����)O��M"E��Ҥ���w�EW��b�&��êtR=8��b<JrК=qI��<	�3qhw�d��v�g�l��uu��;�ɂ��ki{��ͲY��D��m���M��X�Ky���$�_(�x����|%fXۣK�#\xI����;�oRuٹ��jO+�oD�4k�k�W� �,%��
�����RVg֪�m%|��v�V[5J�Q_&��d��n�Md�&�)�F`��0����v��ۂ0a�I��ʧ�
_)j�D��q��.a�-�(��n,;������p���	"�������yر2B��x҅�)��x���5�o?�T9'#�^�x�GQ����`4� qN���&	�L����qo�u�(���8R�9Ǘ1�=�?�:�Yf"��'��VS_�� sv�(���5>�2�b�����e��?
ݣ���!�cna�I�L"���SA�Yk��LMCi|�R~��/Pܵ��J$�+�W a����'�	��'F�k{��Vf��ĉ\��i���Ά���=lv�
1�j&��� �M�H�+�rr��"�bK���v���ρ������O�k�C6��f;_Fr7��F͵b�-�]ߘy>������A�y�Y�\26(�jI��H�J��'�����f��YE�^v�r�`ͫ}��x��n��&B�0-X�~���ui������0nQ�2��x���-~	�ñsQJ��M�I�����X���Cu�*���$M+���m��^��D	��<ϡ
1�8���v�aU �8��{�PǶ���Vt�v׼]����vV�͔i(�C��3-Y�[(ĆU��#�UM�����s����1]L��v9�j�i��.-ɨ�l�d#{Ì'-�+i��-U%8��T��t�8��\V�&�����-�_�~zj��\�4Ik��(c�`�}�P��	��	�Mf{�^���' 
�kUD�����]2P%K�p��ݞ�i�r&�D��U�-���ڟ�����d�D!ʂ��w@uڧ���prb�r�V��U2�	�(T�����K��X�����q?�c��{rezl�6#�zo��5�C�e��u_�|m����$O���$�ZpnG+�j��%GzTR)!k>"�I��S��H�a�	�S����s غv�ƚ,�&�j��h~I���W����-DT�J|���=y��˪�.�F#d�O�
��U�	M��f�g��ss��&�9m<��A0_j�
#�Zpdb2�p%�֚�MUf��y𸍆.����?6��j�e�]�T�
�L؁][�/斺���]�¢=l%W���x,B:��{Y)�,�*?GT�,�+��j��`$@��+���K��Y~(�����~X�:}�+"w����a���\��8b�Gd�#W�QBt�����O��^íW59�7���H{\AU��?ĵ�]v󌬺�/m�5~�u�Qd?]��KP�0���0G[{�M*�+� z�J��F�[3tcMI{e�$�EXR���r�#.a���lË�k�!m[�*i���C��M"׸���&6�����%�{�$��x�I|�-@�S��������9d�p�*E2'z���n\�lT��Ul�N��S��EC9/�g�+T��^L=i]���z/\�X�{�N���!g�*��M��\7�#&&����eEj����Bx�*�}���4�lI�MrꜢSH�U`�ٸ��H��W��\����������i��+�Dxeq3�j=��!��(�H��>u!��(�e"LGe/+��#a6��J}�b|�Lr��'c?h�6-�&`��q�(N��%�6'���-���^b���{�nj<	)d�,�|��t�]�u 	���Y��ݓ���L*�|/}F
ş$�#|G
u>`G���%��)ܩ��'<�E�V�H#�v��VO�X(�0����o��q$�!��\	���h���23�W�p�
��p��H���˜e���z�w�������;?���{�폊�c~V�l��}[��ʍ:>��̠�?��	��J��	����|oX=7��wi�'+p���Jm�V����beQ�͖� G���M_0������SR���c�QbP�����W�c�.&��ٌ���W�O��Zb�R(���<��z{�j��CFR���1�y0���'�}�c��yص0��;��>U�1:�(6S~k�	}6��DPa�	G����D��@>P������Vq&��n�s���)-e��t��e��ga�4{�	1"-����78���
C����:��<�-S9/l3HE��C�?N�bg��vy>K�O5l�bv@丨y���D[��~A��W�ꦭL.�ֹڑE�d���
�Fv���[��2��
ޕPV+�n�<0T)�2��_����:>-���E�m�׋c}�P������R΋Vb
��U
'��NM�:���a��u!�W�H���#s�}�elA�Z���0u���1"M��٪D-[�$�^K#jE�o��g����7Ll
�N����&�x-�&�sz�j�m�`R���[�?�8�`��M�qK<��q�z�Ķz2��J׷�Y)��B{l�ՎZ.r����Nb{�W���"w�{W4��5�"rQP��Y s�D�<���1;�Q���.���n�������:a�0Os�˳��l���VǍ��s�E�-Ԃ\�JL�#_�Z ����,�U9�؂��V���
�I0�6�}戏8�zo޾��etUq���>�+�
C� �1�vKV�O���-�Z��P۶X���9� X�0�H�
Ds�E�����讵��R� ޜ�H�P#����ו�PN�����o�WAЎϵ�UH�<x� B�S=""Pfm����!��|�Y���jPbR	��-��L +�[��:İ�=k��R�`�;����Q�Tc��g�/���r����c����o"��	�����{���!9C��,u�!��G���njz�I���mvX7���s�^x}�LH�I'��;����>F��\0�ݰ�g`j�����:a�4gi�/�c`��>r �2���;�~�d�m�+�nXU��<4��v��g�-���@�hT+�n�"&JGU�����%kl�9����	{��獐�Z�M��TE^T�2�6�YG��s��h�?��)������'x��ȈAOb����Hg@&�����v�N̨a��L���
��-l��G�Q��3�J�N��g���Z�<��nH�c�<
uo�i�����<?��UŇ@F͠M�j:E���s�٣���i��>���}��S����3hhQ�� a%�]��t`Z�>XI�_,((FpW��Ӂ%����̎}��B�<���΋޻�q������'��JoY�!�A�������E�ܳ�}F~�����-�����4Td�#��ܟ�J$�ņs��?�>�Kq��Ԉ�v��ȝ�%��)�-�Z�I�g�}8�чb�jP���0�ؓNS���@Z��U��l��"{�/���X�M��i��ϘZ�"p������Bⶄ��ȴ<����`B�!��F��TT��y�P��!A]>�RG{���p�I��T�8�`ɇҧ2&=�·g����
��?.
���1�m��cR���#�������Qq���dA3te5(������Ҹ��H��@��ջz�sq�<�3���ȴ#�8���	]�eX�Olj�M>��%	�S�E,���LDh8���9� Ct/C��g$�0�o��u��P�fy����N��+��M��&��h����b,ps��l]�E,M�nȟ_�dx��+�{}���^���ͲMU�����	�*�����-�3��,ku2{��h�� ����=�hE�n�p�s�����?��m��Bi	SCۂ)�9tk�"��k�2�5�1_4�BQ�����xe7~M�i��'�(M���F��>����� }��I�455}�'�_�9#��׏�<j�H�*�%����gj�;����h�ANr��K�+��#Ag�')�{���~��K
Gj�R�,�mm�ԡ$�Pʌ=�xו�}�B���M]o��jd�Z�3�C�<��y�͋Br�+r-��V>�q�>E��'Qc7��x]�&!ll�&:�<ЫK��e%woZ�X��ҧ�[.~��ʧPJ)]Q�Z�}��:��UU��ڜ\�Er�����	�s�W5�g�R_=�Y��p���r4�h��S�_;$Ѩ�ngI��@c�ה�A)�D
��{��\��}�OF�xH�[�E��Q�:�_5?���%Q��Ϥ����U������&n���u~�:@&�p�Mu�6�̉{\u������'��� �9x�A�.��lX!rnET^�, `�q�p���^N���P���@�W�s�qC=j7B�I�-&F��"�7�J��,ܙ�4�v��a��JH�|�t�����ebfKL7�� �%��
\6�;;�t{���@������cag��A����B��f����0��0�BDH9{t ��b�F����V˷�w�����|����b�{ۣ]�c��_��F���v�<T�m�o�1�N�r�}����9j\�iz����q�����%13`�yg+��@;���Ylr&- P��Z�1�=p`N&� �!�v�Q��Q�#�	П�t���#��_$,��&n�ym�Go�쩠��;�"�\4k�&��?��h�`׮NZV+�y�#�=��+>l�RO
%�c��+C��u����Τp��;K�H��F�>�S�������]Y�W�1�-��;;��$/�2p�1>��!��R��\x����<�K����6dNM���d=:�K�-����`���5i�D�J����LM�&��d�a�����w	��Q3�A-�|��@7��gy�%X5�_���������24$s�@Xnmપ�ݬ�fPg*���BY�@�sH�O���q�^��fts!{7�i��D�����M�W�m#��N�4�Q��O�6f�a����d�I�3w���B#��}L�b�H������$!([��i�q��?����K�%t����v�t��{� ������Y�D�k��44�5�Gd��Z�^�N�l�F���ù��+B�V�� ��;�'!jJ�@4�1/\/bKf<��;E'j��7b�t]�8��H K2�M<��I͢���K�ul(*���;�=sx��W���h,����8��d������-�'�I����#!����6B����vx�((1b3.R��OX�^#�@�zBƟц{|�BKOj��h�����K�1�����eE�k΋&�	$	�z�P�#S�2�U�lڨO�p[ׄ}�4V� (n����\U��Of� �f� OL���3J�-uZc!&��i.Մ��%(�/�6efԫ|�K���m�7�
�-�I�I�6��Fu����)&1���9"�i����Y=צҭ|h�U�	�������M�hB�$����U\i۝�Up�d��l�b� A.
�b]���~$� �u���ڈo
�M��������FG����\�5��!���e?��v�5���x�O���3Ei�R띬�ݏ� ����P$?�O&V�1�1�L�������+���y$��O��$�X/>gE���R{�^�Q�̀j1��n���A�G9����!1U�EX���{�1�� �n�RΕNy���L�)��(�IVi
G��t�u��v��f)V�E���諊rӭ��,����(�F��wA���/`�9�%d��_!�����$O�_�W�LwH��T��m��aS�"����6g}��e '���t����6���c#,���X �$�ƹ�e �@G��c��[�h��;HX��+��O2����9t?v����l��3�1�}����V[�V""PG"ZzO�\z\X�8aVW;�cֳ�2��5b�/#�$��ح.������[��,��3uH�o�����\x�8�"��π��:�
��@��i�6&x�wO�p4 �
Ū=}��mWh����y���Yt����|?�!dEk�O�!�T����v|Jt3F���u��ob62��A>�1�1K/��9��,7�h>�;y��	�t���s�y�ky#��7۷�����nc�fF>p��B���hY�J]6����"���W-��ы9�o����>�L�UiFE���3���^�!����핓�;q}�t7Ni�chd�W��׃��":�ۤ{|;��k��	M �[��*/�����gu��k��SJ�F_�9ÿ�	����"��ay������l�i��Ku$@ 抗,���4<;����(	G{ڝ�����yPbͭb�Ȉ� ��W�t��W�����Wj���h!A�ixM�/���9�BX����,�HR���ܟ�"�l�/b��2�"!�P%M/��>�Ȋ��Eb�Ynj=_pE�=�#��,.o;��d]Y	�Q`�lꤢ�8�����V��CP$ɦ��;���ϧ�'���_��M��=�׶̝.o�ׄ��M {�L;E�n�ੱH��6�{R=�.�jg�\N:.O��}Ҙ�`G���a/�M�z�V�h,W�Ի�|v.9hT�j��3�}��h�횊:ŝ��2ϸ��e6�;�)'�b��:�j%���σ�E�q�G�V�_��{�A�l��-��w��n{��n�<�qs���-kq��ς��%�y��D�V�:��n	�K ��osf)Ž���`���S#|M��
�H�T������>��ucZ��'�"O��~&e_�����n{����S,�c�9��;IEo@��7N������
c,k{r�_�z��Wi��ɥ�	˶p��P�{K"X"Z~3bD�����$Ҵ%���Y
{N(2��P�~E3~5Z�yH���T[9��g��KY��;���9.�k^Ł�uf�����3UcYt��~��ch����nc��JH�I�2���t��>?9��\��h��o�!�e0�{c��#͖��Yޠ�]��d1�+�x	��.I�@��>b8S���v@ԃ_<��j��$S��XD��{��2�j|�����p��5��.�t�eJ��;_
R�z�2G	l��4e^��)6ʀ�&����S����[��(�� ϰe�������_K�A=Zf}-)D� �am�U��N	S���w�_����7ݖ�Nl�\B�����Q�)���|x��X�R�?��3J7��'�c���R�kMv�_�#�n)�(x�*ȱ�j��!?����	*�������t<�T� �A��~���`Ȉ�״t���8:��yg�-h�tL�H>����$��� ^��m�h��P�;�,��h����p����<��!����a��7�唓@�*�!^wH�� ҥ��������l�,�Y��a���'�	�Yl�n�Xd'�S[�$���_[���$q��?p)�v^c��?�8�>*���4Dq���*&刵��<ZHd'jF9=g;S~jý�b\��g���;l^�pFc�	��!S��q�`�5斿v��#�=�-ئ���F�y�!�O�F�)�,a��qJE�ۤC��>�SQ�UK݅I|2ޣ�FK��è4o���a:��a�1QN0��9��1:.�I��R�P��{>�I} ��eO�܇�7��O���4��0/(�7���~�!�>���ZF^@Gj0�D(ct�s���k�� o����� ɷ���H'ʩT���8��>�y�mvf�}����= L��XQ<*���K���Ǳ�q��j�zF9�Y���u��ɏ�ڹH.{��ؔ���.�9z0��ƚe���Ud�q�=�J,��"�`�|.������;
�/BLz���jhp\���{u�w?7������JJ������ R��s����а��pc[��7���@�ߣ&���h������@|�������^&4��t���B�fR���M��e[.*N�DD�����+g{C����j��?�{�������w4���_��1��=q�;�8\��4}���	\����G�:�ю\�����0��:`~��p,#a�$���	� �x�ƙ� ������T���5���z9�t�,��E�)�]�S�r�=ȗ嗄O4�(`J(�f�j}�G��CO��AٌmV���%q���*�h�jI$G)a��&�rn�D�Y6!L�W�k`G78�[��6��(�^f�1����r��W:�@�̄Oc�	��d������v(�1�J���A\��Sg\�2胻L��������S�N��k��v4:9cE^#��*O?��DpU�����U�:�.;���/C�-�Uv>}¤7�a�KA4<���~�Yՙ�R�%�-����R�N>�森��<�~M�9sXo/y�spT⊜R�W�v�~�u#	�&��yHQ
��P �3��̪e�e{�w+V�hf�&v���wZ]�5�0�]*.����c�Hu�2ʠ���H����+qUמΎ�bN��Σ���C��� �n ���^s2r��K�\]Ρh�<�p��5���4/���ƈC4��heqX`?�Kz�(�+����Y��̉�rG��mo�0��kG����1q}��=�1��7 I�-�{ÿ��� �}��I�<� c<9Ư�2v�]�[��R����'��ڌ��L�`��&�e׌qV̱�uy3q�j����E��|���d(�6^�h=���ҁ:�y{�@�I�@&+�9�k͈�vM�KM-mpX����[G���0<NZ�3~ސUΎ+�H2�K�Osc2�pF�vV2�����9o��+!�F�߱s˴��Y!cZ�^d6��k�e���w+�*�]�w�.U�;H�����+�|������̲^��iK�f+��d-Q��5�����\w�M1��#٤��MTm�X���#�#�ٙrq�a�2D�N���%�AbbT6&���L�U@��3�����C?��}ie�?)�T��$\<��j�%�t��{�t����7䧜eQ�(@�6Y:QB+& i�dzS���
�@J_�A�]`��L�N[Ʀ�-�*<��T�E�-߸t��?"S�uP��@�ls�g�y,�󺖂ߚ 9h���џ���x�ס�F]�'2$�/OfK�����E�+ԙ&C��30��YB�!�K�VCY�v�"K:5�x�̂H�V�O�G_l�6б��n��r{�2ù�8u�Y��!��i�2�/㧀�Gx���/��y��S\U�>�9� ,+����=H�UG'�i����S�
�����P�(d�Zw�ua���;3�����Զ�a3��[����!E*'Z��G�u�����C���[��`��nI] F�Ҋ�>��8߾ER���D
*҂�I��=�FK��z���uTː��y��
��(Y�J��VޏU��P,�Q8�7���6q"�`?����D�xÇ�6os������=� ��G&��L��*y�Vl˞�yAL*?YSG��)���0I?��"X .ǿ�ԓ�0�?e�rj
a��a�<�Z����5�ZS\�7p-y��H3�,���#>T_,6����ov��ZC�M����{J� ���g�D
����:B|�Py��k.{���u٥�Ԟlo�U:5A$*�|_`�QJ�S�nG2(hG�����~�Zm�q��sŒ��<L�U!�o����HSZ�å�|C�'�ߎ��8�O�BҩCé�
�`1)���O:,�}� ���p~E_錐�܊X�!�t�iKJc�ē������������?A�/���P�����&��*�u�OI��-+�z�P����uj��A.ƨ���gS�"c��+�wn��HC�v��c��E���!z zm�t��KP��vC���K�0�P�h����h��L�4�G����젢��'�3�j��ͻ�I"���r��8c��h�����ar��?&c!��U��#g.v�?��t�H�᷍�����ɼ���ԋ�g��ջNCF�Dr�׊Ԑ�B�0͞�����Գ�a�b�8�����e
�|�ԧ@��#�_���e��_K���L�OV8R�Vd�e�z� <#s��2���2hD�DE&���<E�z���Ϧ�M���LԞ2���uw�'F�V�k�-��=�g�X/����+��icWԎ.Pb��N�8�鷗G,3�Hi�
b*I��?s�9=�ڤcB.��b 3��.�heZd�aCS��'Kg��	xqHE�&,(�Zw���&���zɶ�Xt���	��K���T�}�絅��b}�SE�Y����;8r���e:DX��O���z�v�����9_���b��r�g�l��Š<�:����C��d�Oܵ���- �I�Ց��>T#�^F_��O��Z.>���bT����L�BZ��\oo�|}�d,K<wxr/jr]�$�h_�a�_��G���ʄ�w@�w�b�+�`��T�B,����`E��+�MA���:���V����~�;Ҟ�Uq�Ι7	��	��s�4
��@�&�9!qҔ�/۔YC��? KM��]Q������"#v�-Ѯo<�Z/�����F17���d�^�5�z(��o���V �'+"\>�y\�B������H\��w	D�(�,wE�"��J���Wη,=��}\u�슘��<��:;�p�e6Yʇ%�06�L����k�7QH�L�� �I9}]G�r=��"��K���.��'������ZQHK�� .Պ��D���B%����0�L�|�^�DXINq���}���pH64N��d�R�i� �|��ׯ�_+ ��(p�����IV΋�Џ�}
t��K捷I��^�T }���2�^�"
�PX�)>�u/�'.�/��dcS����b��C�b�K}dv�W���Y�6�����u=[ϠO�
דּB�;d�yTI������D]�8i'u=|����)h��۵<b�sy]M/�=��BGv��m��ɦ�3��z�OQ����ˎ��хo��m�m��up�0��o~��鳎��Z�(�#�|0�7�t0�{�b%���wm>�D�a,hN��g.x���Sd<��^9BB�7jF�9<�Zf&����7�p0$�G�^�!���׷ηǉ���#Z�d��(�6s0�'��o�C�|"��4pXs4)��+��,-J-ӈ� i�A�c�f��Q�6 ��)��6V�J?�/� ���u�d�6�������N3��hm��,uX�#'Dj�-�x����#���x������F���GiI������rWɡ �)�/��E�S��W����S��5k�S%����MZ'���.��|[�d�j��r��Jm:n
��Y�E!��~lx�'��I6���dN����וK]z�1��
.-���s B�x�;��q����)]\1��"�΁��EZ����4?e�#��;�M��BR7_k�h�ت�UR>WP��"�t٫��.�+�m�)���u^�l�gP�5ر��E2�T�`Q@\�\1뽷:����:=�8Bl�2�8!n�M�W�uN<��BIQ�<{���oX�s�(!9����M%�Oq%x�������F*��Q�\�c��L��|ѫw�Q�Kbߤ����	�P�\bޖ?.灳���s�Mf��������	��*� <�2>6sS/�a�K�k���;��J�V������D�v���*
;�f�`���߁UOB�+s�-M�Ϡb����'§	O�$���l��Ϋ!h�&�%��R���U���*�?�3P[���a� �c2������e�M �=jw�o��Y5�v%��l���#�S*&v��ݎ�H�<Z�g�@o��n������$�9I�hk4ɡ	�F��m�h66�4�>�d~�n6��)�{��<�Pu�ǈ�/�.#~�<"D	�E�挊���K��R� گ@lS�Y�qhik�"��E�q�؈=Pf�;B��~2�ji�,b��e�)�Q�_��B-���~�|	��`~r��ݮ�aʤ��+�HaΝ��\�)�E*�k�W�u.�x�F�m#?|�Fԗy�ǎ��˳��!�3�K�>Q��Ⱦۘr+`�9��M��F�E�~|Jk�=*��T+��{
z���G8�@���B��|GKi0�L9�$��<��H�#<���֞�7��گ����w����9�NBS�K�t��ᛚ����Fև�^�����������o� �3��ɶ�B�0�r's���-u�_����@u	"��?���m��5����.<��j�2����oh�6ѷ������b}ۖٺ23)HѪ��V��\8�I}K���P���P��y�	����ie�凈X�;�<���a��/��V7����-��EHQ���
k��sP�d<lx	ԯ���.1/mU�.���U.�Q��������]�EōŽ�`/{�`Lng땞߭� �%U�t����K/_f��ݵMW�MLW��U�>	�B���I���4c5�FE��ݸP�2��^�'�esɽ|��W+�QOȇE�Q��MN�L��Z���J������)�,iΞ���q���Ly%�CiGQhh���ӷ�oTuo������0��f�^�(d}�5Yb��#W���5���W�|�Ry��z��&�ᵩQ��Ƒ-7iH$��m�=H�)�Uj�ӏ�G>�7o�bFF?�,G�����o��jn���ԍY��,�ڜM����G�:x�s|y}$+�¯��E&�����2��NG��Ꞩ���ΏZs�7,xR�\��_�W~-4e[xk��D�<�},J�M= �{D�Aěߢ��G���k˗�j4U�&7��B�Ò�%ਹ��|��h�f��3���pD�X���W�ꬃ��q�n\į�z�u�F��i'9�$%��J���Y�� =��k?��
���tU�֦��HL�Խ���_]�&XJ�h?�Q�*f�۹�A��j���3�^��!8w��a6dx1�J��[o`�V�G6�!9�/�g]ujQ�冷�c�x��Ъ٘N=��X�B�b��
`-���-_��{���D��x{��b�η'�@�b�_DV ��Y��O��u')ygW�1��-��y��پ�-���d-K�l��̍��8�s!�ВZ<\x��/�����T]�ȟ	�{@���-=�m��;(��j����=���)�^>O��05 {v�k����&��=�68JAŠ����+���P��0ꕁ�B��8,����l�|��S;H�\�$h��a��jm�1�9���W��G���m1������D]E�U�7<���K4\6��dW��έ����!����GF)�{J��T��`����J�]��Iߵ/|��;�cOߴ{ޒz�R͞B�8��c���l�S���J��)ُ
5(g�{�E��4�TD��	;-"lU���+���Z֔�0�\�Y}�b;�A
Q�R��Y&t�_ÍWd�Y G�baܞ�,C߳=�hQ��T�>�����`�@l��'�N>���L}�4�Q^��3U�܅I\�)_��l�R߲�C3��J߄�dB�T��X!	�����m�y绣�u�;EӀyR1���G0��#�JRh�CN#�to`�^����/#ga�O�������uGsqb�J��П��)]��lU��������U}��ܫ*T9ě�gd�4;�\O������5��}�Q�aG�����yC�����}Bq?8�/�B4���k9n�<U��,�`]�2T6jN��8�:���a �WXd��c�7p�F(ן��L�"�����n��`Фl.���s=��F����,m꼾�S3���ۖ6��W1ei:x�����k��o�<�+�����_�T	Da�&�1�zY?��;��أI���E3rFO~�L2)���q�����-2L{�E�I���$	I���l��Ae+���d��U�1���"�*�������`���`9-P���4{�u���a�T4�a�1�C֙@>�F}�%O^KĤ.\�C������R˸�E�� Ub��R$S�G�Y�2A��oH?ԐuͥKD�[(��<Ҿ� �?���
I��z���?��VA��f���~t��Z+�Q#n/Y((�z��L���_-�/����8�q�t��f.�([�C]�"G]h��vL��mSNUa����f�����D�Y�H��G;�����5t�Z:KM���XNYo��0>)��̡�<f����"��v�E&�}� ��B�3FrC�(�N��l�c��0傴};uM�2��g�j�խ?���k/���-lj�}�n�I���z��/4��$��(�r��%gJ/ث?����4�B/�}�~^n*R%����P���;���}5.�h��zM5�9���!�8��/�2z��6bE��R�AjWP�-�S0�����ֳl:�,u.3j����*>8;n�	=��B�re������N�RL�h�	�ʒ��T]��壉m3k����bg�[+������A/���o��k50��J�G�!��ņ$ɡhz�2����yl�4��0Wk}7닥���T�!�������*FFw���񞈛�eD.C���OɊ���d�������c�S	����8Q����r`�����u�'��F��ڊMC�̑sw��|�������o�V�K)�򦇾�B��g��RKS�������B�PB�j98�Y����]�5�:p��;�Y�kο-�~nm	��ӭ�鳛�O\��z<� o�1T�ۺ$����~�ܝ��]7��V?߆���>�9��&ǋy:}�����t�s#�߶W�n��ug����9x��$�[�����6%o����u���i��y~Ce(���u?iR�_-�6�\-���\zU&<��R���Żډ�0�݆nj޻���-�|���
����jr%a�o^&�9'��t�`�V�N�1F�8�㖣W+�P�H����8�Z꽳N�Qw����`L�����v�M�,��8����Pܥ��dZ��ԝ���d8�:\�h���3�=�D>g�aO�����R�N[�jd���q�m,Ӳ���0ID{���.E9f~��c� ��$����C\� �T]�IZ�b�쳜̦@N�c�WP�=ڵ�G���c�O��6!�b�v��Y&�.�s'��fz��[?M��&���]ߖx��<^,'>626c���H�vu���tHZ����ɗ't���|Hc����p�1�@@r_����M_��v)7�=���{�x����R�]��(΁0鰊�#"�&���n�_`чKF.3�C}��p�t�HCcV�Q�~�-��h�+l�\U��*C]@]E��s/�c�QY�sť;���2���Q�G�T����7����3�}(�nڃ"MʎRsp<{��0��[֐�F��~���Mݡ�E��R8�^�� �jf������7�r�ɹa��M���r��S?<���i�p��������ͳ��@h	����%��@ Z�eQ��P����<��,Z��X�}�s'�c�f9��7�W�7�ƫxƓ��7=�ڙ�ש�k��Qt���'��EB�<Y��;FhT[�(���v|��a4��B4f'�d�av�]i%=웍F�'Z�6��z+γ�d�h�~ /�:��0y�?Z�}���b�Z:ۋ����%2�&��@�𛛟����fe��^5�Ÿ���U9��ɧ���Rqz��;~�O�璉PRL�j���[��Ԑ�dx4�ȳu�� nx{�����e\����?Ȧ�$L1��������qN����iw��||�cP#a��@�+��>�\�l�h��B�/�,�)���J�^�r�s���@�N���wT��x6�J+5����{#���2Ѡ������	���W&{������`r����� �"��${��J���]�Z��dǮ��zKw�����Bp��;��w��0�{�ˀ#�I��.���=P��M�F��OwnV��-�ƅΎ�e��R�z�@M�V��9� �@��T��%$�ucY����O�Z3����2k�d�ߝ��<�'[�-��L���Nxى�����2O�I�Uz
����3�k.`�Qo2�+�����Փ���F�Hʹ
"
�1���yڰ��A(�_�F�"oz3/<��7Y)��ӹ�������.{�3���	�EY�p2�E���K���%ĕX剭�gc��I�	��?ԦY�8͟���"������XLs�Z���֩l��B���p�t���sU�(-M3t���c���l�4�nB=?Λ �>��N��~>��mˑ=<@�H,2�]2m0�	�d߁�9qEDʝ��z0�˪����ܩ7H!O�Q��p@���J���i���RU�$��y{���ą�oaJ�uq��۾���eV,�t^�ɓ�(�]\/�U�>c��ga��	��V9��/@����B�S�ȇ@��:�E����v�� �.����1
�.q�PA��(��6#�C�B"�[y�_c��V��-������	v�mvǭ�K�$F�������&V6������h��@QU���/���:#]:BzE�Թ+Ʉ�,��Q���[p3P�Ćh�T5ʫ�אsV�i����6	�J ��1���x� ף鴷2�����w�QS
gϭ����&��
e-�
��P*�.��mľ���sl�I�&;�d��t�d��s��I� ���k1>�+Ku���_A��m�'��,���~H4�3 ���D�U�b]��C��'�>�+HIT(�\#���9��*a�N�����z"П��5t9�@�f-Ƿ����~ų����)��ꂌ`9M����ආ���칧4��M˅m)O���d�UV`���] [��k@����f��縀�"\o������em�;&�3��|�:R�k���lk抅�Z%ôT<c'�rt�]Ir*G�i��
;�h�ru�
z���ߑQ[ܪ�-���M;�` �x�@""\�qKL:������F�>�Z2���Lc�tr�a��^l/�ONj�I���*�2M#�v/�#r�uM�����#m����R�Í+D��~_�V:5b|K��-��N�,��:w_:�	n\�\,���G?G�४����8�ZL���J�y*=�(#d.+����O�������;�Z���(V�B�T��S��V��	�Ŏ3(E��y�R�v@�������ch�o#\���H+>��$���� nFs���b����o�w�	e=�f��������E� �FW
��Gd�W
��L�>�gL�E�c*|�����������mKث�xm���g[��?9*3)Rp���M�!�v�͵���c�^�*]�� ��qB���:���q�|iD��Qe��8��̘ m�kaa�-��BV���Nha��S�;�s�L�h+rβ������S�C�a{9b�&��
\cHK���?�ܜ�p��&�y��n������x�d��ߎ�.d�،\.�Ƅ&��"��)����7o�Jh:'Z)D���V��is1N���=�:����!cʑ�v���6w�<�m�?�_*q�|M���c�VM�aE��5@�~��W��3��=3�!tUݯ��J@$�&����9E���
M��̩k���z�W)�a��Ɋ�+�:W��Bv� ����[�E��s�b!B�TR��f�	UT<�����b�#}M��&�Ȝ3<�"P}O�������v	����桩3L�Z��#xD���B|X��-F�W�m��<}Ő]�(�s<n�F'IcL%=X�^�N���`?���Y�FWc�S���R���m<?��\Q<'���v�Z:���힡�\�d=�/�Y��W+N֙5ӾW�sVo��T4:�^TlZ�a�ʄ'�1��LO̛#�U��r��OWnQ�y��ò-I��M��b�+(��Ǹ	�/#E6�v�E(��&�^��i�5�Nҷ�}���v5G����㝏��/���NOU�o����Dw����nx6��1p��b�p
/����粐4�0� 4�4.	8�c'�)r�b�볏�Akzj�x��<�XS|��Ι��!�����25�~�n@w����d���)j�Ŧ�I��P�v%�z"#^,�k����K�c=vD� �ҁD�$8b��͜p7p���72-��L��8r*)zl��jĩ���NSh^��(v7�*P'�s}�X�zK��AiG\x�%�w*�YB:r�z�H�%�FzMz��� ��p~ʚB�����@���<���g�z)N�d����u��\ܸ�(0h�a��@��,���O~1���&�E�m���aP �Q�)�͹|I��Fv�P�u}E+$���H��4'�Okp�Nm�x������]����e��[?�	���R�`�����ՌI�ł���d���߽�(���Ah�zt�ZH��Y뎥.N�k$���j*�Fm�\>�'��p<u�Z\Oi�-�����x��wMQ�љH��)>�:B%��H~v�_���TSͦ�ʚV������4���S�k�Iz���,["˷lu���ݓYC�ɚ�tra=0-���GB.���^]c1�n�K  ����Mq\�"W�� 8v���]J$v���\*i�J��/g鶈�D`:bـO� � BõW�NǸ~����"0"���{�C��c�����-����WC�m�� 7]��-�%�͵}1%�=���l��d-9�2��]��|�a�щ10�=��V������=F~��#>�A�Z}����f�ע���6��K`���1��2#s�}�o�\ �XQrՀ]��PZj��U�0�K�	���S��-��!J�̷�O�}��g��	�N����7,ۧ�:��;��m�j�y�@� 5�gUE-Ek��B�m�7u��s�xI���X-W2	WMh�:��.��x�U��AImk��J%�y�X_HX��fSm�@�S-��; �-��Y���p�>����̥�,lC�n:�J}�~����䱅�Fztn���%�����ݡ4y^�8Q��:u��;����6������U��O�J$@^��?u$qY����k��-?�.�M�}֚����V7��)@�Z��.���	;�����mm�.�_��'����雺�E����Ӻ{J��W���c��}�����:�R=M���3�n�m��ßG��$��w3:Z!����� �;���0S�eS��A�H����tr��<����y���EΎ�S�;vU�!���%�͢����O]���RXe*�������=K*���P�	v�a���b��l���P|2WW_1r�ۇ�:!��AXP���,��Yi���2Z]�7�������#�w<���Gv?�&�,�G�����	��@���"+	�t	��,���/C�5h	oJ�n��(����l���7y§���q�f�	�w����T����AW�����+��<V�s8�`XZGޙ.e��4�P�t"]'�-
 �l�y�Z�� �r4#�z��<dzs�ΆV̼��P�Z 3��_qyM��w�Y�P��F2��Y���%��+�|{�]!�Y��{4V��y�̃44a6�wV����: <��;?�"��_FGUz��tp5E���.M�*��݄ YІ�t�y��<��5��MQ�J�P���K������2IXZ8��^�D��%9��넌�T��f�`q�������dr�/:���N�k͡���`���-[tP���[b�%Q%{O�#�)\��i��P5�EeNw�>�q�@~��{%��9�׫���YANg@ׯ��	�g�Y��	 9l��7�H7]��sz����|ji�oܥ��̴��i"%�B��P��s��RLB`��JeID ��_G1Z�'ǧx�lw��h��>�"����,�A����v�8P6�hD/"eۧ�ٰ�F+ك�78��RP�ҭ�=�c�>�q��"����p��om�B�3|d��\e爻���m��x/�HĨYK�M�b�Z�'p���WZ�q|*��FJ������,�$R?�v��g�ৌ�H��s�q��]��ꡛ�q�.�7�e���'�hF)�<Q��Zr	,X����:'qi���[J�V�x:,%������(�	�
�TCx��͈�mL�G��덇���RV0aL�<��r���6�cx��K�=����p7���;���xMXa��_=ZR���ʛ��^�S�>��]����n3���:�Q����ƴ���)�2�_�Nd���C*���w�4V�ɥN꘩΅P6�:[)�����p� ��Q�;��s싫+L���qJf�	�d���ݨ�A�/��\�am��B�@����P<%���NVx�&<q^%��s��r�jԐu��{Z(�kb"�W� �P{��v�-��}�XM��)�[!��y� �6$�ڨíp�`�����8΃�<$r4�!��+�� �GB��,� �r��:~ͫ��-�V��Ɩ�R��{��B�b�u�������ֻ�6�ܳ���-����0"BեYY�{���9'�U��٣��9�5�a�r�����+
��6	�
a&j�/>i�k�]Y����I%u��%XZ{�^�A!��N���Zp�	��6���hVR����#�cLO�ؤ~fт�7%�y��
*	��B��z��?�B[0�(�K�$�����X]�a��J�6G��D��{]Rkm&I���.,���'�#gȞdѳ%/�]k��떚��D�N�+F�a춰0l!��(eB�*Ӷ��n�	��E�v�j�Q���0�����{w
=�dt�[_t�C`��q �Cn�/�"G�����c�
�(�ŏ|�eG�����}���֢ܗ���fϙ7��Y��[haYWN�] h��x�o�6��/�5Q}u��b�\2/��dZ�>��^g*���8c�{�S��x�R���-d�B-Q�, *�A&�]��V�l֘��� Vs�fxc��r�ώ��U6 M�x��OP���P�D�<�`xz�K�)p�*�2w���M�lW^�40����iJb9q�@k�Q=b7U��~Bcx9;ҥ�U�� {eus1ȹ�I��:���7V4�/��W��V�m�xM�Z���L6Z�4�A�۽�>.��Ю�ZM�mA��٫��%a�'9V������)��#P��u{[�T�������M��E���J45l�λ	�)�Q�뙨��/C��.^]��^�D�q��~�WVr���O�[ވ6.�^#KB~� �˕�
�|�1
ŭ�?���HӺ������M��6`��d�L��kq���EW�x�2:E���M�可���������/��:����_�[m��Ɂ����p��5���a�vesn$��c��D%Q3���@l	k?=���I�
�~f�ۄjG�W��q���ô���[���$T�JDN��&�:�����7����G�G"�E�ۦ�E�G�t�=�c,��fD� �7oA lm�ve��I�/�n��9~��A<�Y�axW8�t�Ԡ{�8�O�ܫ4��`B�,2S��K���eL�,����	�g����Vr����D� h��`�w�2g����$��r�]�VX�a����N�#L� L�/����	.��?$i���nsζ�$i��BdD �zI�� ���"��9���0�����c� I����������X.I$��M�o�#i->>ܗ>C�����_��F'4eك,Xow�i턾'��PXM�5�En�����e�p�DQ�O��.���"i����_@���vk;V�Q��gp#0�����-u��tWK*���Z��U��F���Dg���IX�Ц5��圣�k�:Y멄��e���G�^4�����!N�j��G�$����rB��{���}�J���e���t�'(��'�T1 �n������3[�t�����:��Zꨖ�A��������I Y1��XM	�b�,qSLKBh@���T��~l6���\�Ì��n���$�?*��>���Q�3S$�]����'���=5�]���[{}�H�k��:}Ҕʣ��&6N.d��T��ƈ�w V�㄂�f����~i��t�B�����J�{1�����1=%���i�.M�j��0pv�~�"�8)x2�TP��!�A��\�����0�O9Gx纄�o���i��I���&M���:#�6��os C~7W��yVF0�d]o7��jͶ�hn�a �ܻ#�<N_�!�����uP}�z�f	|t����W���KPY�6z=���|8�@f�V���l��՚u�l�ٱ��s�	L�k'�fJ9��r;�Dg;��1s��O���E�^�~��]�(�̬�~����eNt23Y��i�j������-/x:õ|�W��ڧ�U��>%��He�t�`�a8�DL�$rs Gf#l�o�Abz�A�d����o����������ER�Z���"�JD�t�Z^ݡ�L8�`n��Pfk0����R�L{N���pE �L`o+g2h�,����߹m��/�� N��n�\��
{��dT]R�jlu�Ɯ��c���ǌh2c���ǳ�E�W�&�����5�n(�+M�������������{�y�2p�"δtϭ.��I��轡���I�+��HD��,o�n�z�(u���+ܜ����1�d*xI����2�L��G��mAD钗kئ^5���J.Wb���h�s@�jJ�W�h�Ư7��vIY��'��>St��̋�3��a�Qq �;,ö���.��0�NQ
&xf.�:���Y9x]�����+G�X�l)�����U����D��6��H�"�'4�;�C1�^�|�V'��ʷ>˧�\�L/�P)�0�������:Yƒ��~��x��&-�j�(���j��*�I��Y���xT��ilL�o�0�g��:T��Q?�B���	9b�X�W���R$�g�I �6��q.��e��<�#�S���{O������K�\&b�7���%e�'&�-�DAR�q�X�pi����7��|�l��,:����.�����O1H|]��O���R� $
D\��q#!��F&�#���ӡ��_���|�)�V��v�N)`q	��9��ـL�"��X���R_(�W:�NH,���K�Z�,q�j�T`�KR7���	�"1�X�4,h2j?^��P��|�c��b�����4&�����T:=:}��`Xr� �D�� (ZX��<]��Z�����dY��=����"h�ᴽ}��X�^a�6�=�L32O&0����=H��Q�1���z�Y�y��)������j�P[77`M�f�ۂ��d�Ȗ�s�(�Cyrxw�|�h�K؅��X�2LU�h63��Ve������ʒW�,jE��ԙ�ꎝ��	j�����ȣ�֗[b������>��V`�����$�F�S�\�
7y�lv3:.��%>�N���zQ��<{%��G�u�Dy�e��EQb0f&;밠�x�1�3h	�Wq���N�j�@�d}Y2AVv�(�=@y���+~�޵�EJ���H��p�L�Fu|��w�;��i�N7�rY�vD�y��ӊ�*��'��y�����Ӈ�^�:��:��8d>�v�{�1F��(���I�b-q�a&=���F������
]�����R
�^�鱊�q�g���ː��Np���P���hO���wZ�}�+�� �����
1Ԉ�2�t�3�F�+���_m\J��(M�� ��[;p�����!�Z�Bo&/UL�l⌖F/�o�t�(�n�2t��%W�S��)gd�d��L!a����IT��7��2D=�1�,H�%*�Q�������ԒH�Q1�߰J�F��#�� �)��H"�Gֺ�$m  V��L���4���lĵ��B�T�=u����b٦O|�F�YYA��	g��z�oK�%�:� ׻��m�������"�!�GP���u�3	�v0U�˗xJ�_�w��o��Q�����
&�� �tjt��{ղT���⵲�V:Q�Y��txJp_s�9���%����x=j<��7�Bj��<�T�܀�+�a���@p�Ne�d�Դ�����9���k�P,�k��V�����Oh+��&���/�3�򮪃'� c]����=i7���*x*y��Gj�Ų��Ow������x��O�+�S� Ԁ��|�MH������B��1�q�V�c)|ǩI#�
,�!��"և��;�q�_�ΦN3�l�m|N�W%ߜh�
n���[R<ߛ��c5�I���ze=�("c���)�X��?w��"=���EB?4/�]�%�B�D��"_ۗ������y����֛���
CmƑ�g&~���%zhK�!3�I�fDO	�3�����X�m���<�0�(Aw\V���i�(ˇO��]|8����I�,�q�K�e/!�lu�!�m��o�tnv�坲��Աv ��c�E�`&ۖ�J��qd�$Xb�	M�+�i��T 4���X���Ǽ��nt�M�}�&e~3��y�Gb�5F��(�k{���[Y�w����v%nT���J�\���	�.>�F)VTd���ǎ绩� �����؊�&c�q8~�������<I$�NPH�\�i(��#��AQ/�\��{d_x���I�޲�g8��>hf�b�;��s�Gv�l��툝��[��n'���%��|�/�ׂ�G���y[]�f;���k�K^�Uwwr���@� �&�uB�Ґ7�ދa�l#�������,dF5 W��s$�,�@c�Lhe(I�4l ��<K㫧^bש�Q5D��2�Ì�����UHޜfP�tK��. �gb_Q��O$��m;����I��d3�b̷s���\o�
�>ND�b��ƺ�j��5 ��8��n���.n/�B(ϱ��i3��gj��-Sյ�s�j;.�V̯������q+֒,�^�֜�9�������Ċ�e*<~�k�O�9����C��a�42���mm7��� Μ�o:Fk�@\|��l�o�E�y��������ͷ�{�1pv��U�ſs����	����2�F�p��]�����r��E��}r)mη����E8���,��l���Ͽs���g���$z~]I��w[��l������R��-+6O(UE%�P�3�!�����9����l*4y���L�Э�~��Tm5F}V?U���vD�����n���E�ʶ�Łj�b'�*amQ����ƾ���A����x���bV���6�nT��(�YQ#�/�y-��{�Z�i�˷0@�Y'����UG�c4V3"E0��y*�) �/��'k�X���4ђ�D�W��M������h+#�s� �P5`�.��U7Q8�'��ҠαX�a�.������t�*y_�3cd�SV���5�5�ǵYӱY��/��]X��l��Va_�"J�Q���u������#����:9^>��f� ��]��MM�ְu<ez}�D|s��0
̣<pxLH^r���
�0����_;*���N�q��FV�V��X0�5K�{dӧ��p����K�,�v�P����̝���sTw�2��Tn{��NEe�W�ָ3���FdD�6� ����0�}m#��X�{���XB	H�~\;i�0�gP��mS�0�x����~���Aab_��R#hk��@���ӎxY-}9W ���ab�'�xZ��G�FnewjF�V���u��a�M��Jp�?�u~W(�ms��1[p�դ"^r�H6]���`�OS1U��H�?��O�<_ �?��!#e�8/�J�X!��v�12�U���GRc="hx�c&�Uey%�<��֜قa��ݬ�')iV����
m=ͣ����9rS�QBV���I$�c��L�Qv�% <Т'ww:��������&?�8܏sV&��+�j�y ��g��|e���Sqo�B�\�����J]I�H^vR�����:+/Gm4��Wzॠ�2�h�����e&I'|�=�u�S�^A�ܟ�n���=3��G&�Cxݰx;��əl��+�[�ĔF�.w�6y|�C�Z��n�5we�!�O4�q4fe���nz�� ��rQ��CR�h!
5QAPx7Kv>F 㱯��q�qJG�@�������M��9���s��J��j���Xc��"�N՗Cݾ=����2�:T��=��⠒�#��݅�x�ibF�	����[�M[2J�e}6��{
Ua��U����b��Ӳ�J<��h�Pf��s:�{_6��o��k��$u��=?����-4��Q't���b�te�,T�osIU��;�Y�U�ShK���G?�)��Y�I_�	���o�A�D��J.���*ر|Na�d
�_L��x���V�q�҈���Oc�mM���^���?�,yΦˡ��m+���C��O�/�M(�f�����cm�Р|�Y 9���UأQ�fVe�X��v���kX�6p�o8��1���+�N2M������f� JO,L!�)b�ls�X�^Kd�?�����`�Q�bٛ����?�[�$����]���HPx����$~ǀs�8�_a����b}��~��(�	n���!���u(�3x�N��b�5� y���W� ���o+��z�V�q�GH�Y:�Q�&WO(.��\z���DD�Le���uU�d��p�R-��8ݶv���,H*�j̫�Y�9�D��b_�^uO�F邢��偓t���̗��&D\d��5'4&�N8�SN�*IL* }�[7�;b�~'@�K3yI�>���g[�#.�<g�&3��X��[C�1��y�vW �(J���\[XN�1�#L�G
/�Vо��*Гsl[���0X�S�,�T�.��>[��ܒZn|Tg�☇ᶳ`��י�iiH2�M��	(G�)�d�O�R���7�'�|��U����q	᧢��,�����"L��j�K�C�7�g��#r�>���_#��������2��./������q�&����g��_��@�I�k�q?v�I�����{��������<p8jT����N���k�*�d\� (��2���w�y��{�j���w;v�c���<���Lj�0k-Z|
R�j*.M�+;�i�f����΢��d�t�؏V|(5����/�H�%�P�^�y�Ը��(I�^D$��zӬ`�4�ZoB�K�h�Z�������{}y�����;� ���"��_Ds�h^�i��⫂��[�aDX^E���kq"�%�n��@�D��e	F�l���),����`pt����MB�R�O��aM�ġ&�(I��H���yA~��V)w+VʌRN�R��&�'�<����Y1.�p(d��/#������a3~!�Al"��f�/]��g�ٲ�R�J�}�ġ���3���
ie����:	[<�_�����d�>r��0s䱅i��*E�/�nX����;��U�Eb&�^:!gj���#(���
�!PH(WJͭM�b�W�
���A5�cI��zX�rУ�aY������J����'���'��D�![H[-G�	lJd]�c��sO��@���gQ���Y����mţ�����i�CZ�Iz�o	T ��s���y�w ��\&�n��V2�Z~��c{B=�%�K��܍�0"�9�Z���B+��hEV�'jǴ� /�?������y���'�K�/8��y����UtXݥ�އ�g������/��6���^��ˌ��]�'|��}���������j��%ƈ���,��\��0�ѠQ����N%��l�yU�>���A)ZB��`#3�`�-7��M_7����.nժG����r��A�>�"���YА�_�u��z-�{��G�=q��<S\@����O��T���L��	��Y+�p4�]f� IJNI0̗�|�����,�w`���d����_UQ�v����kbK���Q��z�CП�3��C(q0��k�ŲO>�rޠt5�b��^D����Z%�9V�f�!�����q��S7��\\�ܺ5�P@��-D)Y�d�����(&���#S%A�e��Q� ���ԶcOkr�_��?n������3�J8\a� ��bo�}���	֟?��^�K�d�f�+4����Ub��;�T�����"�.qw�űd��Ǟ%�w�փ��� .h����⅒u�8>����4�$�0�[r�:�Ғ�b�yHQfg=wFj=hq�//S��f[汄C`���o/m!7�F0�$%h��m�ϯ�����j{?��ځ|l��Jõ
ǟ��T��&"�G�8�*���3�� �w �[�S�E@��L>i>N�),�UOp��T�(���l��Sa�����'���ђ������ߟE���}Zq䓲����VS<�\#�*Ҩ��7��E�M	[��W0�M�W�K����:9oX�T���8+��[#��tc�^���]|HN�׃�<�b��y*L5ř�k��m���f��e�G��tU�ѿ&�C�B�F��=ZZ�/0���ؖ͡f����<��#�R�v�ػFb&<� ��zu�>�.z�m�4��Uu�y)Nv% V'uW�:��`��F������5���4�ac��;�K>�w	��8`G��BSZ(Zfu����2VoQ�}G���MJ�)�k䅿�W��]Tv��k\���)��aN�GtG>����#�*�f1`2t>��*+����Q|Q6Ě2�$�v����̴�&Ś&�,H����ϝ�/���(=~+"�#�~w��V3�Մ&D�v��u�'��vX��d���K�#s�$��(V������+s��	c�s�� ������1��8�[�o���$�Y&���ܝ�l��3���o�s����4�j��E���q��Ix��z��Ќ����v}��	$��[f�_n�Y~�HP�.��E'�K^u�p?�TAr�1�o Q<=窆����C52g���Nl����`Y�g����
�E���m�z%l�p E���� ǐ-�R����P�P�3��$Ȳ:e>i]�����s�5������i����+�U;÷St����*�]``RQPy�mZ�߱A��@Ƽ�`F�,9�/�F%+�����ޡ�(�%�a_�� ��
k>H��� uUA�(}�^�z����.��LJqK��}�N�ƱZ�l!T˨$�[��0��݆փ�wZӵ��`r9ׁF�s�*�6�iKw�a��ZP��h�t�e�)[�U��.�M��n�l�e��@ϝ|���f�HF(��|%�{�	*�a�=NA�d�x)�W*�AИ�g5ۛ���~r�	R���)v˱�%�C��j4v��"�"f�'V�5��E�����7�Ց��3"�̸��:���q�XʅY���Jo�<8=�;2�����P�Z�d�d�7���\O	�vQ�,=QLz����M����-�&�I�}����Z�P@�pc~�k�[��M��˓�s��Ͻ1z=z��Ի��4?�u�K�%��(%�R���Y7��3��3p�
x�(��|���]8��0^�|ǜF$՚����I\�ouq��a�s�ؒ��E��ʰ 9+'K�o	�)�l
K���9?H������%K��o�L��j��yI񺩕TǽFF���;V���j���-��ݥ��251?[��:|�?�`�h����؆�;�g��=�FS��Ŧ!0ׅ}�ΛL�;�k�;?^6����o���ꨯd	��	t<`U���g����wů��n�p���mM�"�N���p��#VI�k���>
�F z66�=�@N��z���w9'#br��ae��/O��BA�7�ڮf{��c[GLGZyo�[�Hx�P�I����G��g��L*��U,$�-�Z��ѧ��~B�(���@�#VۼK�/:��,[�T�x���Z��=r�<��ԠdI�󙠪��p0\;
9���c�aT��7b(�OM�t
��gM�+lA��Y:Sf��|�41���|~]*q�b�G؃a��Z1�J2!f�A��o|��J�Zc�}<���+[�>�� ˦�!��W>A�其�_�-����O'�*�+���]z���--��01����h��c5RH�׶�\D�!E�3w'���V$��Y���w�2��O�s�W��B��ES�i�q���[�	Ĝq�r��9s�	��Lt�r�Sj��T���?�u�� ��L��^�REv�Ѱ*Z��g7�٠�oa�������C�QS��R���mL�� ���j�.���Ĺ���8Ѯ� |��)Z�!�e�aw�2�/�EP'ك���Ɨ�D2A�����+63����+|����@j�:"ڠ�@��5T���pPjY�Wl�)�r�漷�T��gqMu�`�����J�(f���=�M
����;n]5��]6��K�H򥗈��jJ+i���,�s�*�\Qfex�UC���L`�To�%j�"B�jD*�q����������C�W���3R�f+���鰲���=2�|M4p ���Tu���)�f�o᩼9�����!!��`@������|q������0�#e�!��-I�q&�0�H9KCιb��IlҩHW�#d+�QaW��X�p�n�=Ԣ	63�K�E����SO�/2 ���5�a��z�B�����Rq�d.���Yļ������B�����x�ԝ��5�ͩ��<�H�����@�o�|�n��[��jƯ���i{����	MP�z�8>�x m[�N�ܓuY��ʞ�'҅�[N%S��c�>�+����O	�~�z������x�\��;����S��Ko�)��-���dra왏a��B�?�g:��#-��i�d9[B��!MT�y1��+���ll^�e�.�g%��x��ڸ12C��֏E� ��=j�&�%Ծ0̃R�Q�@?����gǵ(I�@��ί+�;cbfu����6HNS�Q'�����DZ����yo�}l��%�`X���Q�.��&e�9��i7��G��P	�(3JEՈ2���x��N�R���ל?�p��%ߵ�ӄ"����7�9�\~&:.4���T��D��E4�Sy�g:��@,�Z*^��%���;y�@��ɰ7�(m�cq�~6!ārv�y��r���%���4�*�N�I8#)�v����ޟ�y���c���\'�$Y��\�~����p��bm�� �a�����S�GUK�Hda�縞,>��<������ۏ3y+�X���p�bi����� ���;+g��Oϟ�@�O��"�hE�*?�@=h��Itb�:��"S��c�ak�U���1��q(���0 ����`� �|���<	R�@����4�ncܥ����+H�L6W&�fO��y�M�E�]�	�/4�^���3�ϊ�dtR�}	O*���:�Bzr��,5�%�}�uО�Z[��T���h��?9��YWèNW��"hf��Eͱc��"���?ŋҩ�%ޮ�]=�5_a�A��z��BD�I`)!��T���y>���yOs>�%"Q�}��(�<��]�I��%ZH�q<�9]#��H+�C�&Ĉ}�uy)���Z���������W�GO�{�({z�ꔷ�r�xGw����]�Ӡy�-{�s���=�·�7��2��E=$��@6��d�TkN7�X�[DIو���)�+�� _����ǟ�����~J�i'��!~������dD`N�9H	o;}�Ta�n	ǁ@(���?���3vL�ŵ�D#�M�̂�����B��D%w�7��bؙ��#s��%#��Z��ׁz�v���q-���S�?S�p�G@WSYcg����C��=gLy3�?򂳡W��[��i:s�TL�6��D�}�=�����I��������wƶ�� -���Q��FJ�{3e��V�4le���=c�T�����2Wq��yD����Y�����}*�'[Q*�E��G�T,�Z�P���t�Y� ����	��=��HI���朞b���!������Y��@�=&ϰe�'cO��P�>H{	�[K*~Ҽ���zo����3��9*�Zտ nN����ʹ���D�����J�9���k�7"���3RE���ս���WL(d���E{��̞%�R��*�j+�R�QD�D�gO�v�'�L#�JjG���{���yi�_Uđu(V�G++��FPy�͌����[vg��#3�{����Ϙ+�4%��B䮙[�Mq�\�kfv��OsNPF�xYqݝ`,l:�����#;�M��I4Y��0��U�T���k�\[��T�aw�tD$��To����9���%>]3��RQ��N�.'nȞ�/+�:p6+^CE+g��G�yiS�����c��@�M�<��
p6���b�
Y�C�"_��J!�J���%kS����ӽ%<�>1fZ��YJ�,vѕ�sD�&
�.	n֣;�d���x `�3��2>�bZ����V/��R���Y����(���\��n��T�������l z�d��}l6���"+[̽h����W��ܦ����c�����1�I�G��]��Ma�}��H㙽J���y�j���GA�S�����%J�OT���a�����G����$~���B�-l�Vj�� 6Br9+ּ�i�(y�k��/�*Y^��BG�W�Me��e��#C�ļk�������D-��\���E�2�mU�y��=�{>"F�xi'����=�+Y������L)��w�@��B�<R�(�����♚c�_��
j &847���i�˦A�������!ԌJ�^�K��,rR!�Vtjr��+�b�o 3��k����������%��i��BB��ȷ�gT_pds��@��a�㮰e�l�8Q��X��J����Y�o�k^��p��җ�s�z��^P/�9�J��]OtZ�7a�� ��T�B<�i��lF��Z4yM�t��F��S��&[ĹFj !4�6��a��ӵQ����_�R���U�p�L=R ��[����R<0s�
TZ$�w�|ut���cZk�[�=�i�y�&�����-���F��M�&��lˢV�\>�p�&���1����WJJ0��f:9&����^4|>��[]Nsq��_�w�W��E�=� t,��ě���F�ƀ2��9z���oB���+�2ہ` �� ��w;Й�i�Z����<�&8\s�8�_�W��˩���?������1�Y�p*u����D�e9��"v0�<@Ct��vp{��:/�eJAo��{%#KSj�!�����fg�#t�#J����b�u*�4D�����~�m��S�$�`g�;�C��5ڜD�x�� �oY�o���|M?�S}�W��(�lW��{1��a3ȯ�p��NsZ	A�}�漆���񧛯�ɕ���Å����b����=
�؍�Li��YbV��9<�R(x��~��aG�)��4^
C�.�IK�T�3��sG����h��J<�V�l˻E>�ŷ�и&���u�#�@3�Дo�.��$7F�\&wP��*�3�
��<(<�-]�Ü��]K_�"�_s�)#��v�����7��@���%�	Q?�K�92��4��S��&T��(R�y�*����S��E;������<�&��j���<6h�u����w��M�T�?)�1��8�8Z�����` �MmTRCJ���0��"���\�aW(.8F� \닸�3�v8̊[�{�����a=�}u�����烿U
�(��.\�Ǚ���S�?�1��c:�W=���4U�eW���@��-���F�ȷ*s؃���PP����6���Q��Qd4�\݃�\hLݔ�R��2���	bh�o��o��OYOx˻��uK�՘ޫ��3�~�㻨EEh��n����yg&��xb��3�v�O�QH(<!���Ze���N�h/�`�i1�6��S�5��Z�󟮴'�ǽT���G HI����b��)q�_�-M�Q�oXhy�[Ý�[�@�'���]�����'
��������?>�V��U5���@%N*F�r�˵CC���$E/$��ȉ�K뮭T��	"C�_5�Uٹ���/8�',hq��^�����Y����M�'Q�"�	�X�-uzъ�-B8<H_W�¦P,�u������ī�A��'���ܮ}"�11�&��v�8��Nd��|6dŠ'�*�rV�J�t��<8V5���+�d�T��C9o��V���G����`֭c�F���6%!>�d�)��G_�#x�!�զT�����)�s9Q��=�q�{H㇒$��{�fG�윍�n�OI��.Oi���#A�!��pEڊ�#tz��������߀m<d��hT�����y��+1���%y׍7V�Yl~��T�j;��V��ť�<�ӞU�`��0����na��b���S�w������V^�N=�S�l��p�.��D��,�E��"��_��I7����%*󌋗�����([n�(�����h��&�G���Rc3�����M��M�e���w(0��!E���ՠ�O]��%����s��W1����p���I\#Q!åZ�6K��F:�6�#��L���v����O�`Y��4���@�غ�a��2*�I P+�6� �O�b�&a���E��ea�w��f������i�ݮ��H��y�H��VZ\2k�m����RЭ#���]g�Հ�ln����E+�e�%r`x�]�szړ���0�N8�������==q�o�)&4|�m�`k΃�~��'�[���Fu�*����g̠�56���:���ޭ�.H��u+7V0�Q8P�ԯQ�t^������t`������G�@ֿ_9���2n<���]�f�=)��.L�Ùox���z�Z�]M�ހ�T +�kC��Sq�F����� ����7���-���-��V���B��:�f"v=���2�1F~�dfa��5��*3�"�ڨ�(�;j��a�z�J���=�Ӣl���l�Ք}~S4hK	�u-�%;q#�	S��
N��/pF�7w�-Q�W5d�#�t'���м<�tV�I"vXN�	���q��=��b�.�y�c����Z�e��~�r$�8f��1���'T�1g�fɅƆ��`�kt�E�D��7���!� !C��ǧ��1�8���4C�+��P����VQ'M'^��؅mo���Mb 1@��0b�+��������\��"wRo�5��D=��Ϥ�0�<t��{qQ�/�����u���p+��)/�jcǽ�`0����Xwz�J�%TL��ў���˾H�KTe��?����}�gB�j�/=	eҫ��WiJ�������*�o�Nޣ�@�	�Rʦ�����w��Ԧq��n;�r]��:���F��~�X�HQ\�7��	����Y�b��,�mv��p<�*�.�^f�`W�3�i:����<l|��|�(+W+R��z���3*�Mh���2d���� ;���֐}CH���c#�:�W�S�lvi1�j��*�Mb���V!��h���{�����4�M�KJx�)*ˀ�O����|�"�:��A��:��I\�AG�: �kΜ�'kj��vb���> ���YU���x�O1�{�D�v�;�����[y�d��V���)-qY�|���W��	�"d�"c8d�m�T�R<=zۣ��|_�D,R�~�̓����>4s���+r�����=���� Q���hQYo3��NV����
��T��':�e<˙(l��\���69��t�"I�S���Q�~��.�G��P���A��b&Iߞ��u�,v@�<F������ƀ��gl>�'�l�J��'��,_������` W��S�O;S�2/�Jp�g8q�<�����'��#Y����e�����G^�~��)M	�C.�X�suJb��銮6qO��o=�F�ZB�m;B�2$�nk��i�4jw���K���d�;�m�94��ȭ碎e5�#-;AW��`n�}Ҋa����,o��ǖ�{���r%{�U������H�$#�������u�(��o�.�9�ضa��1���^X8ٰ�(k�K�VTD�X��8��K�������B����2M�,x�u/� E�ã�n'���~�oI�k3V�i����+g�~����a?�ᦇdc�d^tH������U��ͮ\=C�3#�t��oMp~[�Vx"�2��RH�@Y�U�/G�}�L���Lq#�wo��-m'��EJ�-�6�yɁ��v��iw%q1�D�e�䂴�	�-�*K���]�s6ހ��8�WC/�����	*�"Ǿ��wq��B��t�6�hm�_H�X�L"��T��z��:}7<YX��W���#����t�B���(�������(Ӿ�	S�)�ø��-�@5+��/�&�Q]{q�-�� �X6 a+�r.�ZYyO|�\�"F]@���_%eq����>ȋ7�[�����M��"s�9QY�5Fn!8������v�	e&m|i�:6���.[�k�%C���Mv�K蕙ߗ�gcVX��͍�s�r�6��蜿\�wq2anqh��2���I�O�x,��t"���L`.Xf}g1�4���9{�</��Dj����p�C7��ܰ���9�+�u�>���voϗ�KZ�(���gXI�K+�P|�V[�wi�|lt�u��9H���h:N��1T����s��.z�J�J�p��ۑ��K�M�L��!�ʹ���&�fS��@p~����k )�_�$�B>��w9�"������)��1��m(.%U|��WҪ*SE����[I�H�0��c���0��H�O!��}��m<R�)��c�a�k��7�e}:�����>1j��!F�����].���\sX�)י���av��|W�rw�ձ���X�(5Z��i��:��yQ�r������[L��k�s�SVXxܸ�|2+wp��$m>2�bF���0j�����8w	��<h�;ZϴW��z�4�o��0v�i��O�u��D���stsmKS�f��iޟ�%����S���\^ Du�@E*�ؗ���{�� E�D�T\|"�K��;/"I����y�R�l�3��;�2��_5�W]�^+	���Yg��ڐ�����)�V���jx�4Q���mԲ��W-~(�8+�������]E���J#�C]�=��ѣ#�/"��c�S���1!��fM8�y�z�Ձ�V_�����˦@@�{脴-e'��oC-���soq��ֻ�!��ܕ���]ǊyE &i`�f�s3��
��Rz��ո�:EX�]r�MB����w��#epM��t�n�jesچ�����(�،$c
��s�q�~���>$������Ct�x��e��^Vy�r	��Nk���̩�����}�(�:|؈�a��'���`K��,�V����X�ޮ�^iC:W*]s�nǘM93vC�{� [����_?[&�������%��M�tȃ0x���ײ�~�)6���^��v�;&͇Pr�O�$5�+���0�u�!U��G��H����Ye��F��vU�4�	&�_t'����tAb��R<@�UUJ޵<ʤb�K� �;?�6~ �Kc'δ��� ����|xs3QڷR2_'Ip<q�(�.6n��$o���0s=����ߩ��gD��c+�amQ�_WL	%�زy|Q��ʣ'���|�<��i�(���Yf�C���q�C���~� ��K���Gȹ��h��p���z) ��P�[M��?�w�:�>7\�T'	wv=�0��Ϯ���P�6�`����چa��gE[�<��AWG�4<�ԥG���ɞ���v�!�XL������}ʬE���w��U�V>�Z.�QI\e�\W}�M�3h���y>�8�휌�33��M��.�G��`�^��@���d2�����f���E:/( w,�@"�*%8Қo%�ۻ=�<i���h�N(��kå�M.U�܀0�H���vqx�����sfn�{l�V��TŹ����0K�ݮG�+9�vs��[�Qz��G�.�횴c�PC.�K���ݵ�=;:@i@^�Fa�[n���Nn2�w�mجٙc�#B�]J���f4�ō'ѡ�%�~Ŧ(|�Y�ĖG�Ց>F���Ap�dw������Z=�{F덊�T�S�a� 3(	���$(��� ��HR��z�V(ތʌ̧Q��y��ߨ_V�hڗ��D7Fu����Y��O:������.�)���[�ޑ^4��B�!���DaC��BUs^��^�'��Ğ��O�8i-�a�}v�DW�F�1Mc���*|����t�%�(g"6h;�0��0�E{
Iy�\b�j������z��Eb��c8gckA6���d���ۊ/��l��$K�N��tŮ�c�0_���fn����*���t?U�U�6�JP�IzA�+���9�=Hp� 0}�����f1�/� G�l�-@�p�~G��'��a����F����2Cd���C|#�t���5`�qn�'��|2��% B?W���Ҭ�ؐfWb�� �H��l�E��G���x\�
+��RN�-�c�a�	tA��Mp^Q��l*"C��}b�e%�Z�s@y��,D=Gׇ��!�B[�^|���elW:;��u���`Z�Z�AΑ�q
l.?���&��?F �ƻc�E�&�Ś��5���>:ǮL�g�ve�@'�J��բh�L$wr�)�ĵВNt9 ��9��S���8ҋd�NK��[$�li���L��/DrH9r�{6!�'�����
��̆��c�cz<��v�ҲJ�-O�*"�hiM���BR��{:���~1�#~:`�%gē��s�U�;K��#�s�	Ӯ�����&�^4��(�֦�/���T:�2�mh�ef}4ձ|"��CWB2t&~͕�'Ys��ґ����*�)��K��'�q�n)�=Y�{��I=��[T�ĺ\ς*�EB�A�1;�r��j���ġ��&��h?��,!!��]��j�&"�L�P�=Jr�~*^>��Q�!G��6�P��"s�	������v���]�l�������-��8;X5�9�G�����\���5~v/2�Y���Af���h�x$�ʢb$�"���w�ND�r�lf����XJ�hx^$Q��:9a�R���Rcz�����e�����q��?��j�R���UoY�����eY&]�]ƙG����K��}�Wz NY��/��R�f�M��ꓲ��?�N��{ެ�6P��\�OGW��lێS��UEa��3�����@��G"�Ȼ0���!Ew�1�ܿ��rK�F!P\�+��
�1�|	�}�[��V���d��V76;���GA9�s ����ç�ت���V��e>y�`����� "eox��Q����6��6��@n-ݍ��Vy_ǝ����5y2�H�co���Us��d����4�r���}�5X�}^��'�ӱ̦E�?6#j�vz�xL�O�:[f>�d�2������N��D�u������;1_Y�!vߪ��2ESn}�J,�6��`��v����}g��1�n$�Ol��1�M���[T-��]�I���Ӷ�~��K�X�&�h(EV�x���A</-���@���;�����'e�$~����?�n�z��n�u�O|����>-4j�xsN���Y22����bY�C���������3Z�T�ͺ�r���<~B��yՕ_�Oݡ��$5��i��f���N\��%]�k�ǿ+�!HL�P�v�*cK�l��t��_�6�°!�K94���a���w�<Ȕ1�d~ށ�C�nMu�~�ݩ�"�����Fx-�9L)�۸��|�V��tQ3��J��G#c�:B�bq[��\���̰���!3p�[X/f���y�o��l6�������������]�7#.���S)�)M�X�w�'���T�H+i?��b5�A3��ߥ��������ʎ\6V��PJ�rN8W��i��%ppl�����\��V}�`��[�P���2/;�+�P�3���HA�.X~� a�y4n	�k���:�ݘ�1�l=�+�� !�5���c������עF��Q@zT
�M)?,�������,Q�b}<6�IcX�4��Y|۾�A�6p��,����[^�N+��3>&)��LR�����Gv7�� �y�d���?z���~���C�I�����_	C�=ޙmd#J�V�zuW<
��Gj���0�a��@���Y�N����X>Z�v�@ҠK���b����C�iD*�5>7�*�Hn,�x}E� C���%d$�Y��z� �<P>�����a(�Hr'�j����ʊ�%SZ��&��6�k��rm}}��9�����.)0��%D�\����l�$�
�l5�M/k�oqj��l�F�� `L����W0��ׯcS5O)��$�	�k�྅&�s�|�mb���P��3��R/�X��j��x���`'��h%�o��e�ŏ��$��؀�/Z���A�j�Э�ꊀ>��`�j�����ց`�K{8��sU�����n��V�p~���в��#��:��Ӕ�M���*1�ޜ3W�]|�e��.c�j���T������-��~5��_� XIo�-�D���Y�&5Od"���-AG��j4Pxj�V�xg2�j�6?�o�U�9tΛ�����K��	#a(���%���_���:y�$��%_pQ�|mk'S���[�?z��
��N������E`���sp����f��\)�ގ3�7�~��)�*L?A�9?�=��Η��"v��̐�X�)�l�I����A��U 2ZAA
P墒lӆ�@�������U�EM;.�M����,�hH��6>�"U�Xwo*�3PM��ISH&)��0�z���?�,��՝�$x~�.�l|�y��oOH�rjB��P�YC�`��v@�O�W��B�h/��%)�4a�_^�z�:C�U�y�O��Ⰴaݢ��u����zSl�L�@>�{��܏|����V�{-����y�.1^W<�����	��x	X?�)�7
?�������˨�$��e�`j�^�`y�vJ}��id%f�_�8�fkG4��[r] %9��6�U"�_�3���Q���8ؒ��
�g�u��iU��I7�����PB����P����5����-��\�魽���/'%G���r����ŬHH��(���n���P�D�QVs��ÍZ<�(��Jֺ5�mL��W�H��R�V����)�=�g�a+���I"ˉZ_�se����<�F�� H�ˈ�6�,,8�86��2�&^���5�$B�Y���A~2�xv�&p�_�y�}5�L���r�tnw, �<�~y��C S���ϐ*�d��Oi-W�s�mk��x ���s�NM���Ӵz:��ϯ�r[-��u���sRcKc�0#x,�A�������jV;=��oE���'�T%s�+ߐ�}�U3ɟ�.s~ۛ����]^	j&%���b܈Gy�z.�;mӗ�T9�4�*l޴'�rx<�X��{���U����R8�yJ4&=�W��|�ter�aydV.ݳHa�W���𢕃K��I�T�;d   �a�Ē
^幏��@Wa����>��4m��N�X�����m� �fqh#Ec �J�~a>8���먔���n�D��1F��]�}��_D֯=Ha������I������ip^�� �w�[@��$���Vx�ߖf޴h���k�����C%UR,������/�7d�������lN�I����(��o�br��S�B�nn�f
� �i�\7n�9x�}#���K���f�!L(B�3��T��9	:������~:Zɩޙ���xRt��.��B�4e��i�i5Կb�8������c��j���OE�栬s�Bd�A��O��D,nQh��r��ԞJ��#�H���%��UP&�u���Ldx;���<ӓ+�&&ˉU��a�Q��P�O�á��/�@�`R�R�&���Һ�/�����?6��u�o�r1�,��9��Y�Go�ӱ�)�Z?�U�_��������KFЉ]�\��~	��x?B�n�~�H`��ĝ�;`M�s��0<˼9x��[�rH�&������Վ�K*ҟ�8O9��d�)p��|�s����zd���X!%����\���6Ed)�bg���~G���oQ��H��qa������s��&���%���.Ah�D�G-����+���/�MY�/���e�w��ֵW7��Y�Zl'·�CN�K�Py��� �0)iD���i#@$��6���C��94X/����M������"�P�Űo5�D���n�i]{i��b���ܪ:��4Z7�B�����O��t�j�햹w7Y/Ψ���|���Vkc���w�R�CM�n2IW5Z1\��
p�1�-�%Ӻ
QP�5����̣�Oo�����`��-47� �r� �P=bLQ�jT��Z㺙�pw6zr&�n�:�Ы1�LJ�&���é�a�N�ߢ(���yxqk�s�$�m�H%z���]���]em��X�w��<��ox)8�����4 ������[�]'\�#�����D�H���3ŝ�;�.4���j�*U��8�5��������9<0�8��b�m܂Pb�b�J�ol��q�^�j��dH�^n�X;3�s|YS�Ո4T�4�"8_����Fh��zE-�F�P
���~za�z����?�(��8˰Ӭ�Q~vx,����Ԥ���$5b 12�0���y �uw�/�����M���DWf�t�Ŷ�|� ��ؒ\3�����щN�`MAr_Z�E�IH�M����uUJ����evP}��-�0��䅢��Q9���:�w����`lӮ� 6�>��Ba%y�۟�o��T!U#��I��|��"�Ѧ
(N��Tz �P*ޣ�cG�~ܓЊ�Jq+\�<���}�۫�waw�]tk(���䑺,�4idx��u#J.rYv�xʞ�ul���U�ֽq%��#	�EqC�ޤ������;��!��|,u��=~F�4�vfz5�

L��\P��RdK��
�Ë�N��o`��|5��c�v����'������䂳wi����"{{Zg倵St�d�e'#�[��ex)�[��d%�8���&�7�SO|>�$������+>Jߵ�q��T�z7av�B�{�76{w�i���do��V��^��1L�s�2R�5�}P�v+U������a�O�������p:��{<�l�@���=�A�#Rk�䨇��]�4Q����p<'P��-8���(M|l`��Ztd�HͱĘ	E���R'�9����zn��?@+�ST�?�aB4����w����1�T�����8i}2���"��&���~���������'���_�#�e`���w��\!����ח�����'� F�y�Q������Nd4�>�H�������L"l�7%%u ��Gc	rk�D��%��"5����0�$`��L�Ɠ*��)a2�i�{ݪ�����/ܦ�������\���F�
ڴI�3n��R��Oƕ��]on�����b ��@�����#����F���e9F����F���=���섫����W~N}/t��,��Q삦'�!���?�B�],��{���태�ó⌯ZgP�Ռ��S��zu�j��zKi���8�������0lq �[�g��ލ[�K������H=��ʎ�Pա����s,���P���a�?E#r�l�N��'�Z��0*�@O�#�YҪ%6��{w�/�余��,�TOU��Y���u�5�Lr�y��������7s�ȃ<��
��zwjot��S�Y�U�����n��>}�2_��zt����>"�Gi�}�Xޮ�CT2�;�����N5?nN��
�O�K�^����0*{3��$����L�.]B7�Gs��,f���F^����ۚT���_c�4�*���o]��O-�1��Z��Bu]��}��}��_Mٸ�)>Ɩ ހ�+����-5���1�eQ��RC���9\��-�*�M'u��Qz��I�E�\,���ߙ~[��e���+6��1H��� �������	}�<�P^��R��R>f�d��5��r	�SD��/�ќ;a�r98��yO7��q:�OHi<��)n��r�l�p�@z�p��.-2�0�3�9���m�T���p���m(���YN�͂�;���Qb!�Ǟ� �!�:)P˕�H��-�S����ʏ`�&։�4SY���x.�l���-eN8y6���o~-QiBRm2��l���q�h��f�ɑ�q~NS]���+Ex����;(q.�t� ��2�z��遗��A[�C��	���3ǋ���߷&�W�x�H%fϽ�.�U�ug��>Վ`'Q�a�����U�<{���`#P�B���u�w7*���l�,�,�}%U�l�
��N�,��}M�]�;�Wʀ�o��]�-
O�����<���Ʈ�nr-��*�[�9Sa>P�"Q��X7=��7D�����J*pS���x���s-�Jm8��KV�w'�8E�|v�Ya�5�������f����)?�'�|L���n#�C���'�/|l��f���	l�3��1i�8a)��zG����}��}�y)�(A�1T�O�2;�ձ	;�&:���_h�T�
�O�4�E�������x��r|��,��z�7۲n��+2���r�@.�7����m*[',cM���ٝ��קkx��$�A����_|�ī�\�n��ZGS��W�0E���=�b��H4#Ѵ�k�%V��h>�=X��P��u!-ݸ�$6�%C��=����1�y<j`!%���9�IY������ˈ@?1���!�3����T���ح�B�=Ǧ}m�L.�%0��"i�����gD	�ff��j�?�@E�8[��<�.�˿���yt�֟Oh��X;��H]W>�kL�9�H����D����1���%��;�%�o���(5rd��lIul�+�i߄������=_�����J�՞;�d�'@��:o�K�?U"=��Qa���T��M��.�v=�r�H�c�e��~�ۈz���+�[K��AyQ
u�<��
P�a� �3�v�=/�v&��g�g�9���d��S�g�g��[[���!=H,��j�b���� �Ô�*���4�F��i��?�W6�ID�|�?
��o�U	����+�P�Q���<jd��T?[0�_�|��~�j�Ʈ�l�#%�"�v��۹��P�O�%y���^0Jo ��^����%�=+�AS8�@��cJZn6X��9��#%r���dä���(QZ���_e, �9-�_��U)%�>��P s��R�и�a�f��'�t�E5���˟��m����O*�.��4g!ا+��Ul��M�ؑ��N����Q�!�X�߭h�p�%�j�2�ؠ�<�0ү�!�oH�UK�Sx�L0��P�����%UL�'�;����oJ�p���ZB��OMVpn]�� �i�J�9"O��Ь�;���m��1��ĭ��q�aWO��G͢P�C��c�ے]0d�RE�C��j�V������]��R{-�2�k�%5��9�=>��/Tj�ѰSD�	ձ9�ټN�u���M�C�n�#UQC��R�ݖcOڌS��/��'��:��B�򓼧I2Wm��w@��M2�zOGAM�g㳍/�TC�U��$9"���v�#����H����x3�wU��O�`�b� �[�5�BǏ��Yb�fS��
�n<?<�p�����Z{�yƄ��ԂO�B��2�@(~x,��D�;%�j%�d��z��0�:�+�=!�h�o0��t���M~�+L�T�P�se��𿛹 {Lt�eՒ0�_����~eFT���*��"������<s�]x��������q�x�re�G}}�yB�����L��D�D�C�Lt����X�m�����+�7)񁵫�,�y�<���D�!���RZb��c�t2��j��w��	﹒x�*�`Z�<1A�S=����۾L�����39��G��Z��W��E�(Z{ߘ]@�3�
���y�lC��E�Lɕ���brX�}�-_;�*}s�ׅAs M�˻7��Q�c9\c� =��p�Ui=_�{��0J��*��@�{Pz�W��t�Ԡe�k��Aģ����=�����:�?�h�-�� J�|��o��!5N�bG�Q>���:j��'��7w��s����$T(�����/ɑ�;K�����5յ2 S�� ��]8m?Doo\J�I��5\�g�-s�8����W@��&�
� <�#��$���PD8�E���|@Sߘ��R�,-ЈI�Vr������4��Җ:��-��A�J�L0*�y4���L8�%�r4�E��\^�2^��׋3i.��0���G����;3(�72�۝ɆL���ѫ�9J��sC�ގK]��9���.�C�1�N߁��0�C��	e�.�Ci�e�̈^sF���'���	�{S�;?(���̄F�
L�l�<	���`퀿����	��f���W��rAP9)BVm+Ͱ-fo�i��L/�Ç���Iʖwvo������5��Q��Kpŕ���7�<�^�"�/q��$z��ڃ�\��fy�e�����a+�uO��4�J�YZ~��.������Es��_>붤����]�*휈#�����������y�?Lkw~��h�&���,�S{���`,.
)��r}��q>��5/ӂ��.������
��=sŢ'��"�v�a[m�k�:%�6O�4f4~Ih�J�����7�c�bQX�D��0�B`n
�$�S$�=8i���p�մ�Ňw@�xI�n���`�C�)z�i���_��]	�"H��ɯF�Pt�h��	�x��%��&�7�8͊�n�k�q�h�-�K���_H�2^@��<����#�ngW�#�)���p�瀐���|�+
ES�;�3?��+���Q�>��N~���FU3��L(���!\f@����j�~���>�qqχ�C�C��SK}
���Q�q�A�E4����!�wu�.ƨ��֖������8s�c���h��������q`��o��xqg��,ۆ�!~`Kz�Z��Ir�@f�5��$����OfV������P�q��נ�]�."���L��8�
ߊ���J[lS��3a�(�����@_�0�Oq_h�����Cw��_��9���ѻ�i5��05�{?׭X�)������=rم~E941�JTO4{���,Zh��]�x���'����&�B���c��o�q]y i�"��o��u`�f3[�M�����[�	�8�v��,���������K�̱;�H�1߾^�4��7�=i=p9��x�i\yt/(����AʏN��m����f�zw�b�0m��Y��"�;E�f�ӻV�zB���R�'��������r�B���Tݧ0k(�/�_�~{@a����T��Vs�#]i<Z_���ww*2
�#�h(8u�V��K$\��N�,{��[��j��7�?��&�	īw��$�R��Aw4�ȽH9՘ߠ37����E�Y),aS�ȋa�5�ۻ��6p�,��6�"_u�9N/��dN�I�*�ig()�ݧ�s�p�%4����z��vG�7�z�Ĭ)�S��bŃ��)����Z�O��_PM�"� aF�	�#![�����.u5�e�,)j#�L�3�y�T��PkF*��@�a)J=&���zT�?���]����>2�B�]h[�wʞ+�n�5��6ϰA��Z�Y���J]��q��u����!O �ѾR*?��m��W���ϴ㣻c��v�6���s�D��Hp���Y_�h��q�8������*F��/�.�|Q�`}	 �!����n�?t��GNaR�j�����<�F3��m�x���1*K=7�ǵ.�W�,9���je'F��WE�,�� ��Ċ2SwR�XݨN1g&H�2j+&���Mi�
^�	7�.$�wRu���ʧ����%x���������a6me���y�9�埸lM)km¥<�M���6���1�bp�
�[![��KW�)����N��V��ɣ�P,��zwJ�l�T�޶�M��"ޟ!?�ʛh�E��s��b����_7�Xҭg��]rS��T����X��L��r�j#F�
���]ť~�+��1�g�s���)�
�}�9������3v���[�t���;�0i�}y�$�rh�|�)(%�V�)��^����7�R�F e���ڧ����C� �`��V.)�uB F���:��ܺ�y��%�g��k�m�?�����:�o��FA��j��.�v��;.�S.�D�|��T�
�i�~�,�閯1��逃��Y6��;+��N+��=�]n�Ŧw��vxn`�a�V1k���: �{�[1j
�T4��j��� �pڶ*�T����uQ‬L�=���=�CAX¹G9�ɂ�3�XW���7���7����YčH+`��hdB<��~�|��q�Wɳ�)|W
Q��,�p��02��T��Aҵ�T��_�ALj�	��aJ��1<�e*~PZH��'�"�g�E��Sä�-�5\Y�� �s��HB�ח�N�ڒ��pTrD�����Y�~R|}d1�4CQi4���K ��7E��5t��x��P@���x+��������E1���3�:����b�����/'%�S{���O�I����}O�	��y��kJ�@T�V�U�<��a:���a"J����_�-2���j�7�7�T� ��E�3�n0 ՞\��T�A2c�ҏd��+컶�0���m��v��2���q�J�G����֌L�p-^��3��VU�Hn��pq���^��l/���t�d^���gN�"�m�v�6l�ۗ�gR�r:���*�a�"�P.P���9�<��~
�1�����(E<�����t��[k:�lC�����q����ws�#/Z(�J�,b�3_�ܯ�^�U0
!��)N���W��B"zN�/��5y�[��/�ww:W���R>��c$�S���S�))7܂[ �DV���4������-Wy�JЛUE�y^}�h���q��s�݋>������I�b���\2��G��==�0��A�]+Uu&�������*m��K>fy'?�uU�ީ��*��o�:�ʔF���;�ёY`������F����ie �
pqZ�t��G�D�l8j`L�F�B�.��i�dC讌l��A�K�����H�x�6?���2�>T���N̴ܢNU�J�R6҄�@o�lQ]�P�|�������8��	�/	<�u8U�q��Utv�P1�T�"	���<Z'Vސ83f�4����G�oZ��qW�S��y7������϶�|剶��#���Tj��M>	_�V��Ș�z�ͨ�e�X���4�,�����z��u��RF�WJz�6��<���Bu6Z!�D�s�Fw2���Qz)�!�j�-��R���� �D�韑�D��Ԕ��N�������J��4?���~�H3�XM�����ll���ۨ���hx34M����v��@��i���s��P��i��]��~�Â���El_U̪�����hxS��h�X#n�8W�! $�K(R��D�++�͗��{��c��u�n/�W�>}�_`�W�_�hX�0�����&}&�0[<���-A�
����l���09��ǌ5�F$b�Aa\�����m���(�����	O��e�w*�%_V�'���I�������2�f��	jWI�%Q��mك�mb7:H�����d��h9#��.���M�&�&z���@ !>�����8� �X���
_wѤ|�OF!��V���M{_+���6P����0����«�6���O���A�ѯT�te�oǵ�k�+T|�q�H6�0��U���z����y�m9�6��3�6�k���e30d1C��!"V�oӯ!y�V�E�-Ia����wx���a�3��j��yK{2��!V�`�B:u��p�<fIa!�x�:V~�)z�p�ʨ^�Av�V�|�x�x����:���r8�F�jԏ6����6s��Wȃ�	���Д�fG)fۥ��  �3�p���:�x�َ������@ݏ���C���#�����B����=0��N�j�1;��i���^�s�n��#A�'�H����t\��󺶣Ss �"@]u=�ׯ5�a��B��CEiv0gل�����3R�/�Ws\�����D��Lx<�V�vX��o���ڬ�z���d
��sEf�g�U�2]�{�0|D�"
��X��+�Ý�����d������z�5�l�Xs��V��s���VJr0��ܕ�n�Q�4lҮ��l0�]�@c�R�g������;���a�> �±�(?x�ژ�|�:�y�*�F!�B���V5t�|��tB�]�P}��.N�QNpXh!����bҍa�~ṕ(���LW���e���u�T�)�qo��˸T<�F��0/�M.�#ΌV ����l�8sǢ�%������.ih�X��Y+p)t��W?f��Ի;��+Нm]�����hq��z��NM�?����[���:W<�UF��EM�b8?�|���̭�e�5<��ϙ��"Qn/�jB!$J����ыRL��P'n�	�q��U������<�>��vW	65��޶�T�)SZ݈h�D ����a�C�c����y�MI�o�pnH����=����iC��J�U�6A ۽�}HI�%b����-B����Mc�H嫠��E4���p)s�3�m����&��`�Bj�-����� v�M�;��N���l�ęK�ai�<�Y������&�+��?避\�G�Q�^��v�G1?�׬��Y�Fo��t���i�Kk��{��:c���p�>�_�
���̽��P3xAZ �~�� H*s��_��ef��_�r�#%bº�F>�m���Y��Q٨bˍ������ �ƭ� �e' m~&�
#|ij�ȶ5̒������Eu��1"ᇪ�HR	t�J��#�lGƨc����q5��-��_!9�V�Dx9k��������uRY��|�ӊGBH5��C�����:��<�^��G�L�iR��YG�������6�t�$���h��X��p���U*/J�}u3����:���,ڄn��X��3���p������S�U��YZ�g���#W{�£[�s��p�����,�L���SmC�7�J�5vX�&� ��f��JH����BX͢#\=����_�ƾӢ	��2��
x=�i0E_N�j��&K*뇭��[Y`a$����&���q�Ύ��ـ)�l���N�"ǘjۙW������� F/b�6*����/��yZ�9�A����>�>ɂt<��ML`ԕ��Y�d��
{=��qn�)R�WP�;����Ih�pR�R��a=T��'c���ģ{3k�zM�hnޗ%���1ƶl&��2��a���c���+�������C_��#�
���Ob;��_D�y_���?"W*F̳���������j�g5�D���F3r�Z>k���yA�˵�vo������_����L�ao]�f�j�z���/�au�F�нv�$h]4��׎B�.��G[�[�*�?R`y
5{�~���تĮ��
���6�xbt��#]no7
[�J�6U��<LT���OВ�X�T͠kk)�/aؗ����GF{[�,���z=Mߊ���fsNP��cA��r"�9�����'�c���4�¶8F2�s�N�q�s<��_#{�
`�
&�!�E0t&�k_fÌ��n��}ޕ��}�J��������M�Ÿ�J�ރJ��R��gP�jē��YY�;L��%��=�^��<L] [�����n��f����2` ��2�3K�%�ɹ�̽�~(~�e����Wop�~�� 0��7�+<]��9�pM�����#�ӌ�s�k;{�OUx?U�`!Q�����	�(�`��5�t��n2у�p;��m�B3�B�4���u�8�$��,�w_io��~6��ʙ��׽�(�+gD�i��4u}i��
a��h��p�&�ue���,[<�Q�]��VY��P�����١��b�4�'F��C�V�*�3�v�0RU�Z�{�����8���ȉ ��;a��-�'t��4�cxB�U��B�I�k&� ᄷ>�{�7j/���EUJ�k*cNPH���¯5�����]d���v��^�΋�57���þ��T3K8�i$�{&���J����1aL �&i�ǼeZ���(���7�ؑlf�����m���*+�G�������Wi�gJhcl�� �Ǚ��Ֆ{�3<3^�Υ,ͧfq���I�{M����u��A�⇲C�v�'5�t��
K��Wn��sP���S���9���}w.�{ε.Z8��R7M6�Bێ�fcx$P`����t~��J&!���2{z,W5<�&�N�ugR���Y��k�kzX�[���i�&���}Q\�9��jE��������;��NXK�B�<bh����������&l�r�
�ϗ�Wc��E�`@�P��`o�j ',�ʺ�u�ABn�rm��j3��&���ӽE�Ɠ��d
���v��d�^�5�)���C|��)�R�3��۫z��f�>��a%�W:��]+��̧>.	��
��VTe#s�ao��*O�4�f�P#�錃�~/�
���TY�¹���'@���~1hK���P�6N��֫����QN�P�q�R����癁�D[8��.Ycs����o�Q��
���8�QM��K��7ve�/�>KO�ڪ}�o����=/�9��"��"���o�[���)[�7x�H�<��\��-����m��� ���2Axc�uc��1��3�'�0��hX�c".GV"����a>B:���E)Ov��a���KN1H��u3�ɕ��v��!������_�^͞g��a�Ҷ�.s ��e��d��I�����Za�����M�g���it�W���5�B��૤1����D�A`�:'Z�A#�0��V�Ĩ�)U�ɽ�Dз���8< ݛ�E��jM�B]O8�T��;��@K|�*����W��0JS�� ��5c�O��jN�#_�&�Ta���t��@�;)��g��jFC<*BQ.Z��9���>���w�Cq�W�g����+�f�s6����Zn�V�������Ed(~b�wZ������Qt�Ŵ��u�%޶�������NG�sdk���%�(��=��hMT��w�#��j�'�T�7���ֲIg�
Z-Vn8���D�-V�|�c5Zs&�_�Y�,��V$���{��=�M!�o�3�����f!p�B����� ��&CD3��k�v�^����[ΑZ��]�㍦��(��d��|tԺ��?�񼨖�IM)��V�������޺{�e�(�/W_-�ts�	�b�l-(�MB�:.�ޖZH���9���{�b͚5� @��Bo�ώj�m�Aܽ����J;�F���N#�M�#�����u�Y��6�?���"۷��Bж�ab�����{C�Э+���D@Hf����:.�S'�0omj�9�1��=A-��E�S����u��{��F�-z�H]-��j*����$)uf?�1Y���8HY4�	}�Y�U&����X�/'����zY\WH�M	%��]P%�T�}��:K#@.�� eWN��+7�V�!�!�F5��cS���ѼW�A�����9')�>�M���uL����h�n���Vp�2O��7��������f�Q�uh�޹��0
a��*��LO2�~Q��[:*��f��H����<�ԗ�?-�{y;gY���=��ߕبl�s��%�f��{[��G����^�`��G��*����'�pvWh�u��"� ܋����<��_Jup����寂�,"�ze�
�ͣ����Н�$ᄦIQ�����q�.�q��
�gS	"ׄ1�颁�����`v?�e�o�+�K1����S$q� ��<�2���T�� �Jw��9��#�����nJ�S[e�2\y�>�g�WNV���{��=�\�B赥��R���yW�0� 	�Zv[t�����0�.�<���ųM���ّp����X��/�k�Ok�ò٧"�~0����q��ik���i�"���1�Z'������)V+�����;8�wc�G�HM�EW+6�|�Z�������m��+�����Z[Z`��񎋕"����i4�d���&`p��yD����Z�LWTPm2r��y&�k�>(@�|��h�R�PMD�l����(
{2--�B�#��׿4?���<��J��x3���4>�"���q�fk��CN�Mi��:]l��U��D�t��e<PK�>�3�x���ĚCO�ќ��[��l-�_�;���հ�����;����LEM��Bg�M�� �p�3�Qj{cI�BA�C&?�l�,�ږ��a�m�(�}]��`���qtG����#�2{ş,�Pa�� cŋ0�i���@x�I�+vB�<4t�� ~��0$��v#�D����|O;+��/1��u���PC����ƕ�/�C�v�O��:0��Jy��T��~WHKJ/��R9첱.j��_3�wJ-�q}	����
G϶�Ԭ���]�>���y��+��aֳ�,+ݩ�R#`�(�f�u^N��@��dg��"�%
��2�7ko� 
`�/���kb�g�*T�H�Q"�B+��Ie�eP�7$��vO�$!����K���K��x��OL&rP�0����0H�l��ԏ�M?]��B]�f�r�K��#+e�m@��h�ayyB�0oܠ����5����8�y�t�x �ơ�����*��kVJ���u��� �{* !�@��L	�WԴ:�H^�2i�J-Kbϛ�Nt�����e�jY�4�э��ȕl�����l=��"Q������WP*����r�<���!�R�1��	�+mBU͔څ[ �:�<��c "Ƹ����걂Kp<C̞�#)�h�^��\��֭�0\PAC�F�6�
�"`�/a*2G�5]�0b�k�ϑcG�����	W���|j=��a�ȴ_���?_̥�k��.�z"�L i���;<�ց6�P��K��|U�<�m�ǯئ����s��Ԉ�ۗ:���X�E["M�]�iy��i��.At�?ѵ�5�I�?�i�MBѝWu��T,����=>j�,�����-C��Z���j[�7rok^p��2��_i�m@/a��4ʎ -L���F�-���i�Q�l�����O�v)����o'XV�Yz;���@wQ�oś?����TO'�\f{3��¿��.�<;xX�d�Ҙ��z�J!��nQ\
 �H"-9�ˣ�ٛ=�5��"�~��2��/c�?��z
����wi:��h=;�q=�2����d`c_��$�㙁��q2���0G�&��1�"D�els�vY.�\޷���#���Q7��1*2�][|���ʯ�AA�X{������5���U��@W�.��nb�/B�<�K��~6|~6��a�t�b�4w�+��i^
گ���~��$e��K��E�+� K�TQ
wh�'�E5m��Gu���\�������'��� ��0lE��&Q ��d�׌;�z��$�m',Yi�z������Cm{����p�H�Stj�2�sz['�M�\'&9d/���~].�I��/�CH�OVMUJ���E�������td7
�5i����Vge�;��8@IL�|*3�#_"�<�>�I,�-zd�z%�~�zY�G�O��y$����~�ϥ��Gx,���1�gޝ��&}L�����jQ�o�[(�2z���kxh����;|��{��<i8}�}a�㓠5=r���Q��A���?�uKk�(�p�0r�設#�����������E]d���0�r�Or��y���,�`bg��,��i�5�ssr����zDx�Ԕ�*�$�~�P�7{�ܡk,�<	�r�ysow(��z *�OgP1��.�
Jߊ���g�5M#�B+]K�Ul�j��y�
�����_�\%�y*U����w�L?�i]1#����̢d�P�p^H�H܌�m^a�FA�G��s����d�7�"��JnL�8%M��>�	�ʜ�o9`�O�+�G$�>:��(a+�v�Mtz��	����@J��N��O!'��޷pI��(�[]��%�1?�b+ 5��_�"V�\hPN�0�EC-�Zzl���6��=���'c�ƭ�N��M4P���"�V�S�M(U��C�{�HT�mf[鑯���G�Y�D{G�����Ǩ����5�%�x�K�0ȯ�'���Gr8�&'�"��K���UvT=��vo�'?�P�+�P5���'�G~��1�;�=�ۧ��Q�����ƅE���3Y���*���o�+ i���^���-N�d*�Q.�	).`��{�y���{�꺿6��Vu*�*���L�ƚ��M�����E$�Ё&�2om��Zf��F�R�x��[T���̯v�3D���P��:f4�����F��C�h�����5����Y5H�;=	���r(m03h��^O�ke�c��Y�dcO��WQ����H�(��֬� j��&q�
d�m�J�_�^�Q
�g�0�N t�iuwдQ�`� �Q����	��zn�[���Ǒ����~.��~=`Q����vgN�f��,��&E���(�Ǒ�O��Z��ɤ�N�܀XM���pB�X�$�5��0iЮ�
�Ön$G
��zN�L8��h�z���'�,��[���녇�m��c�{���a����w����Q�o�� I��<�<�a(�g����������!>�_K(�.�VV��֓�I+(�1���;ݱ�l���[(t1����9���/#+�����B���@��+�y �Ti`�5�^��F�M�+ ��`#ꐤʴ�����d���-�	�z�V���N��Ө��C�!�ҭ�s��LVK�x���ޒ�']i[D�g�i}�hdSڥ�H�/�uy����H�=��O^�CC0ѼUen�A-����PI��	`]�� َ���xK�o<v���&�x�7��`���c�����Ur11ܶ�<�+c%����9`�㡢����	Ad�%�p%���{�u��n�t"i����@u|�sV�֫��~�^G=���!��ɞԐ!�@j޿��g�bNbgU��V篽9��F�~�l=����� Xر��������i�^ʺ	�֠ڐٞ�.3Ctj����Bn:+�����7琈ꆙ+�I������rH�-H\K����oa�a�K/yĲ��y�gP��Q]y��!@u��R��R>��*�қ�6�2&CՃ��������{xӹ�]1ߙ;��u�s�0�M��NF}��1ٙU7��6b;����P�v�i��A<��#����L�WS��V�l�KPݞ����ϙM�t����In]�Ĥ f\nK���1�?��fI�Ǽ���=pSdf�s�)�i������Y��'s#�P����ݿ�P�P���r��y��S*B9El��Oz�R�4��Ul���&M�f����^,���Û
�k@���.�W$��N[�
��t]S���]�$]axcAb�8�� '3����y�3�Fe������)�=���K<#\�5g�ꚂR�O�����c[ˣ��J!��y�BdJ��bR��=�nօ}�o���S����#A�8���"+��'�O�]ޡL�ê�7��h�8�)��B\��pT�>�^_��ݡ�����4b�Qa���f8SHH%�d�Z���ĉ���;�~�}� m��lU��rY?��Ӕ`E-�q{���7�1q~��C�Jm��>�J�_nRpk��)�� ->bc�'E�G�>R;��T�=�3u�|����ħ��;a����EA���zSGǉ����j�*��IQ�iz>��*?(���ݺn�if	�k<�u��Ck�l��&��݀%u��Л���
	B��?���Ns� Tk�� �]
�|�'��A
��,j��e�)�q�1���a=؈Vy�~��~
�2U|�U-Jf%�ȥ�Ca��P��EC��Z/�{k��us$��b3(��c��z�pr��(�T=3L�"��Y۴��^��(I�(7�T�;t]�-v�,)��eKSz�>]�8�� E/y���l��t�u�LGߕ'3���̫<U�3���hs� iZ�6�H"�����0J����9vG<��E}D�J�Q�=t�=�R�_��P.�d�M���Z�ѳ<�%�����h�O̡���JR�jH�k���G6��6׹Bgv��7�ʙ�Lo��'�%���qO��x�f5�e���ؔKS����Jj�ka�	ƎO�Ed���v���z)��`��IH~7	S\��{����W 9t@[49�Z��Ś��[,�6�Z�"�適�U����z�����+���S�p5:����Z��H<\�)ӐhA�
ie�6�-ɮR��QV��������8'C�+����\������V��������La3	xG�e�Vj��DhAe, T�Ʈ{F�XP��e�� 1�;�.�rU�4u�!NEYi<�ʂU�QV	�7+�Z�[����y��H�*���P��s`��G}��)zj�wۊ����Tv�99�T���:�H�9�O={�.�@�qH�%0���Ł��O���%�M9�V��f^s�/q��^��T��;KL��C�!<�f/����=j� �]�n����Jk7�$���fؚqL�솎����������� �0�IoSE
�m�k�Z`(�D��ul*$Q!m�.iQ���tQ�ł<b���>����'{=� ��˅���s/�����9��i�s4W'�K㓚4�n��!�wY���;���$b����:.bl�g{�l?tUgm5�"-'BD	rοw�2���e�h�9ޕv��Jej����f9�,1�8��6�R+`�Pr�f��t%F�0��t,���W�]uQÍ��x�p�P��%)���!�C�������%>��go�~����He_����dJ�(��^x�gmMAZ�]�k ���V�����>��/���h[�2�*j�%N�@Z����҇R 8�l�Ϣu�|���p�L;�&F�䁌㣹d'�y��i���#ҵ�/@k�xK���(M�W)L#=�m	{|�1�%�J�6&	��~�˧��L)�2���>��5ϕn��)��.f���� �2�8�f�����֑@�W���R|�a���hUǺϏ8���[���O��[e��+�w��FG�]��s0��TB�Xr|����v^��3\�Xy�:쩢���+ҧZh���rED8?[�����"E�o`������^=��`��Yؖx�F�J:�pr�BR����7�F�P0�հ��MOS�w��	�_m�ё���j��E��T�_ @>�m�x�$h�S�<����lT����Y
�T8b��R����a���i��i��j~���W^C��H8Td�N��80�q��n�LmV��I��Br��r��-B�gI�%$4Z�qT�E����,�ȾXC��IOc��
�z�Jԥac�������{�E�O���"��:�״��`5�3<Lq%T?-S����I��ʎ�,��آ�/�u�~��6e4UycG�Q�"u��!d K+��*Gr���]��W�lM��y�m�Si�3�	��W���4���°�ۙ�����z}s�W�!� �uٵ !�1c �!���k����C�g2=�6>Cu���]Dy2������2*��i&g�p�pj���ࠎ����+�nv�9xK￈����L0�?��p�;���H�ؒǂX����f�O����f]+9���Jb3��d�O[V�=/{k�x�X,{��SL�Z"g��f������f�ǌ
���'+���Z%`g(�g��t���;��8�� Μ����9�;>�-ZG�J������n�ɛ�|�.M�%��o���x�:_FWk(O����01+�E����N�?s�L;���k� pXb�^�ֿ��Wp��m�$�dd��˔t���u/8�m���X�j�j����b�'������v	�[�~��xy�|ǟw�͵J��K����;���r53�LoE�q���ƛ/�QIрf�`�~)����ix� ��m���Ҟ[��-1JN������%���@U"��-�l^�;���K��I#�̹���F�5S��)T9���hQ`z#� *���pi��,i�X�4��ÞD�Ņ�m�L(�M�:7���_aM��$.�_ M�LSz����N0��f�n��<�4T䨤�_J�/G��"5�� Y��a���b�`g� H,�nA�$�铬|�jT��T���n�����y�� ��WYQ�t��X�Yx�W;�*���;���s;fN���u�� 5��vn���F8=ͳ�F��^�?��Vl���Hw������e��u��g\�D��"����:�{cmьt��L0"�j�K�o��6�D֓�"#辕� �����6�������Ð�CuW&��7գ�Z�Pi�4��������0��5�ee�y�f��" �FԹ)7{�M�Xf�?tn�/I�޲V�QT,��b�X�c��nUnI��f:x�x��R���nX�����.�j�J������E(�{�����A��x󠯓'h�D��!����:7�;��d)Bkߜ�/�{c"��R��!��|� �O0$8_�z`@B�Q{���R�m,�����(L@e�������p]0���=�PU��|	��֖ݣ�����b�[� ���&4��h�w��]����Fu�'������hp����g]/u��N'(e���v���M�� �@���LȐ�Z�sd���3�_R�
EC?4�j�i,>�,y�Ѣ%�}��}����K{>_����$0������q's�++u����!�(C�s��>P:=\/��6͗���t+���������HrP$"�}�l�.��<s�0H������Ca^����d��I^<�������O�[���q�;�:T���ך�(2ڮ��70�8�y�ѺqqS(��ᠬ�R�i�!�(\*��Ux�)�V#x�K��&e9�NY�����sr�^Ht�&���2>`[m
�vm^��_x�A@ pw�	�g7����}� d$�����P�����RM`T��~�H�E���g[=/������ԼH�d!�3Asb��k��(A������fH�΂�H�%�+I���OL�<s��i��@*�TBX[����V;�]u[��j�����WjO�m��9!w��frn���F��f�����a�?C���M�
g|!�6�)]O�"2�(R���쳎^�|�̸M#Mr�XO�>��M0�`Aϻ�Ѷ\Z0u7����)��}��A3��l���0r��Uܯ-�k��xT��%W���X2���#9
�#�g��m�Ab�H��t+�++tڲn���>^�۰td��j�ᰏ�Bf��K%)b���tUҊi���b�	������9��K��&��1����k<Lm��D^Yf	z��1��ؒ���u�a�YתR�{�� B�#��-a���B��9 �p���v��g3��n��=���W ���LZb��B�e��T�� sy����GP�'��>�����}'&g�k3FX�'v��=�|=��ϠA�g����cl�iL�bv��z�b�ǣ60e��d�m����v��;�WJ����e���SMf�>�{����?��0���W�>߈���^X$)�9�2H �?.��|�ՠ~��ݖ�=�|�T��-���L�����'�d��s��e���fkל����� M��^z� ٺ�͘��������i���dԑF��-���.��,��6+���9G���kц��?��\k��ti���%���]��~�V�k�]���*�C�����S�c���r�A��8v�1ݩ�;�}�t�����3�0��& lTݣ�3G���и��і2H�?'��� b��1��:Ce���.��{iA��)*���j�{�K�Sg�ٔ/M�*���m�~*���2�C8bE�;_Q��v�XHT�b5���/��Ҩ6�t�߃��Ӡ[37v�s�wל�?��6�^z�c���^=�?��T�X��:{C�_����Z�KV|3}��L�!4�Z�+���$`I���	Z?�!m�!�V>����3A��c�:"u�Qd��Zf�3?,�ϑ��g�v\��:�Py�[���g�9 ��kg�.?=
���'���KкC>�7R)a'�"��E��ӧ�P��#�}D�!Z���>��,^��'�y*�d<��Wj��FJ�V���F�9�����囬��z�Þ2�M1��e/x��R\���X�����/Q�O�)VW�a*��L�CU��v���:�R(�Mȣ"�P�}�~ҁd�����y:ھeR��4�����|��4`QY�yu�lj�ëH�|35
�:�J���<����ݽhM
Rzc�$�M����dB��O�������n���g�f�eܒU�֮���'CÕT>�C���Ӯw܎���]j�$g4l��o ���|iG_��{�3�Co�h����Ts7�35��{:^�l���]>}��r���	�z�6�"�2�����H���g���/40�9���Y묮զ����KL$��Z�1`��c���/�ܣ ��L?��6-��#i0뼿�p~\6m9 Ȁ�dwN�!ȅ=�ޒq@�Hꍤ.7��	�j�Si�ș�2C}���`�E/�j� �}�o���Gg�W�
a]�anb�%���-ڍ'���Vk�~�������R (V��.�Ѱ�w����E2|_�Db �WH� ��r���e��&Z�pʓ9W����s͹�drY���N���AJ��"��1��VP���T���?�A&���~'I�� �i�ٳ���N5�\?ǟڒ/�S����lr������"�`�n4P��%�ΰ���q�w:V�<�G
_�}e:)Ǜ-\Iy�{T��� � ��)�u�rE��b�$KM݂U��*���R������ �T� X�{<�zt�"���-ֲQŢ�M�L�l���0�>t>s;ܙ$_E�O�^�}����7�e/�`OI;��T8.V�%��5n���[뉟ʒ�Q2~\��ϱ���>��B�D��8aN����`Z@�%d��E��v��ӻ���-�mm &k%>h*:��S	�\nݝ�.���XK5��r��,g�kg�w�4��d6�I��	�v�<�N�=��↉����	�'��l��:�h�WN$c$�x��>�)d�	�&�&�a$#�,�{�U_��E|��h�Ȼ
%7���{J(KL�6V���<����=mk��=�V|~��  F1*>�v�>"0�b�l;4��T�k���l��:)ĮE�Wխ�9}����{��؉@���:�����J�ޏ���ϫu����S\
R'`��0�0<yс��$���7�"ݪ%�E0蠺�YQr.+y�<�>�܆X~I�7t)b�nOD��>c�1ו2�a,�_X�F� `�	%��<�T��6�8���ܒҍ�1�Jυ馛Õ��S-U��^� T,g�~T��&q ���*=C�����w���� 7{v#�-|�����֜�!L�:��,��n��jjz�%����S�?xǁ7y��	*&��J� �~`WAEG�����>%f�ѥ��<
q��BD��)���\(pmd�r���̝o�c*��&v��Xz�K�Đ��V�R��
6"������������rUJ��n��["h`�G�<_;9��DVώ|�e5�goal�Nz�%k~�a���@���qMi����m�5�e��8ې3춻�a��l�?�Ղ ������E�Y�� C�}�b�Ӆ�7V�-|)����v��+����m��K'��6�"�V�aAĶ"˻G�Tĉ^hcÒ!���4�o��<�+*rv��NDQ������5��Ӏ4������h�J0�َ>����>��f��j[u�<*�C���F��p3�� ���ɔ���e����C+{�����/H_� 0W��-���7L�p	<L[���=��*
��*C�HG�7@M/���r��p��WW�'�._�S���,����m�;��yU����ij����o�A_�N~���	��)�j�0���N9�5������w�go
�ǁ	����>��&T�5v��j&���V��Xe4DcN��å�ޚ�� 2���延��O.�2(�BP�!�� �n��0���՝�mx�W�TH琞(5�p]Q�XhS!�d�=-_�
���s��A�A�s��]��R�w<����'���+�G����`�++)뺕�/�A�)qp&7p@f��Ɏ_gK�3�r�/*��r�-��q�7ϖ�rp*������(!_��wO���u�	*7H����<���bW�������ي��QC�<%���iw ���Ǡ��u�0	:&�܈�h�N���%�B%���-����芝�uw`�i'�_�oYR��:��%P�i�,x�dm�ٱ4�.�1i�Q�����DdC[B�l���z揨�v*V�x�N �T��/5�B_U(�u�� ƞ�c���e�ǪLMM�φ�i�I��t�m�v#�
 >Tu>���I�b 2|�*SZ!��Ǎs�+���i���ǽd��/�׏w���j=��A��=� ����0�3Wu���m�/l���A˩m��%�Y�<��" '�?Ʒ��+J� J�&o��3VSsoCs-`�)�)j���,�d�1|ꞷ��Ew����ILL��!�$��a�ๅ��|"nZ��N���G�� ̇A�f�g�8��,��.�Q&�d���p�f��5��T�0�^Fk{�h�  �U��*
�$A�z"z3m� V���Wӫ!�k�����@H���0~�Pt62�f�yvϟ֞�V/��۪��!��䷑���/"O9B��zSRp�c��Ѭ}h�i�35������`�*K�`G�?��+a�������yؾ��"d�����Yw)_#�&��j�N��9�GZ����o�Q�	�2�v�E�mo���3
������y��|m,�;~�,���#|;V'�AD�xY���A �(�t���Yk�`Z�ϋ�W[t���Bi����ȅPD��5��7� �ܩ�v�h�,�t�M,W����Ļo�-FrFj��X����
�%�؈|q!�i"��ւ3@��r�=�kw�pa1FD�x sҬ�F�� ���7ӹڒ��� 	�6���f���t���Cm�g0OvA��r$�H��1���r�p���sknN��ʊ6����<��ڕx\G(��}҅C@ܺ%?��x������WEc�d5��ma�ᠮ]J-�z�Ћ�קH��{I��5�����$7���������|9M$��k�<����|K��
ȳ�+�Rd��7�>��%���o�B�G�W!g��4_��ol��Я�wY|�?nSB%��	T��d+τ#����b�9�{':d/ݚ�z
l��玉���}���\�Hp�hy�*|�O�v]����� X�5\��t"�ϥV��%%��la����H�T���~��?�������x��wرO�9��̓[��<��f�s3wGb�ߕ�>#Vx�X�2m�[^�7����e��ٯ'�jJ_�`2���m��!��U���3��dsX��cC\gMy%�^t�'"9R�h}����F@� ���w�"sMo������aDj�B}�ie�34��9�RWmؗ�RL�	��ts�m���+�1����ܱ�p�P0��(�g��"�"'��`�T���/��<�h���K�˂=���_I�}V͎M"Gm��[*R��~ù\��@&����}�0��>�����DS�.�Ɋ��!�yj%?Brs���֯^�d �;�8}f�Kb��ka����V�ې�#��к������vN<�

@�[�B��e�'s��e�W�7EȚn�����a��{!����|P����P�~:NL�P������flo��_NH�F�A*r���n��͙�}yhvޡQ���_ �����üχ,O���M�E�;�bv������Bè��"e�1�=/%��e�0���[�W�����5���Ðſ����H�"P����eQ�ob�yEº~� ��u�;P^d"��=�K��p����zM�b��?�yb�4����(�D\�|���8�炑� �YV��HѢ �����,`/.}(��1�a����R�ЊoS�N�H��������:�NYʐ��Ht�+��r�t�9�!��)�t�xA ������s?	��rŁ`�	f?��,�����*�cn����7��
�~�D��*H�\��]����INs�5 � �O��#�H��գ N8��ϟ<(q��|/�9�g�nԺ_9��Wsi�܌��'�w� �B�*���?��,�i�#!P7���+H�_KI�K�8�
s��QA�ZE���pP-U�d�!,��7��1�;)�R�DNQ �~�ʥB�,`��C�٘�pp'>!�#�B}��TD���c�/0n�XI�=cЊ�`@q�%|sR�}�Ɵ*
܌(���h���fcAG0}�OCZɥ��nj2V0Bw~�K�) ��\��8XUh�]]To"�uetg�C��3w�&�V�ZL�&Ķ6�"V-=�p2�lD��ѱ�~�ԶE1
�R�3U?�/hN���Z7�T�R����\6Y6Di���M�@�)0����]��.8�ߊF�YD���*�bا����Ѫ|��c���e�����d�9���������@|�25 �����)�F(�.��+z���0�:�����7�ki�_}��GE��@�¦LӦ︾W�t^{�S8Q|�m�~�N)ƞ��y���� [�c�s�;��f�Wg����5\m��P� �㍜WQ�ѱ�ߴ�y�f�zQK��\o�W)��n�W���4=���1u��㩞�CLba|��]��H(Z����u�kkLp�����8���m��ُ�S Gɔ��`#��rthp,U���䢦�	�M-B���� �Ց��� ¿͘B�	\qk��B�xp��*�q<�+i���8����/��n6m�~�d�~��9AfTU��R���Աmi�m��֤�j����	`WQf���� ��u�����܋I�ݻ�l&�s���qY�)�Ϩ��1Z�=x-�4\5m����e��r�D����Q5���vG��Q��T���0/�8�R�o|�)(vH��"r�荴A�h��^�dH6>����>�u�B�͞���Dq�i� z�j��$;��8�#Nٌό��z���Y�P����HiY��(�bG�b��t��M���c��O�(���-a>յ���Yh[)0V`������h�o��C�.n��2~���k�ˀ/�6���`�XbK{�ݶV�@����o��l�J`eA��T�)ua����a`z����4�.P��,[��4¯����yp34I�����\ݝ|:�?V��y������ �]�y��ν�:�B]W�]�Ƅ*���m���Leu�]a" �K�sNS�3F�/	b�[i�/#�N�_�2n�`�}������U~��-� KI)���cR�BF~޸1$����;��Ќ]�ɠgf
܉P�E澆�g;�gL��l�����W��/2�˹uo��
�����]ˍ	��x\
�ӻ; �HK$]UX�Ԍ��\M�6cM�h��1|�����2�F��q��w�K"y1?t��K�z��~'Jx���P�K�����U��)CC/��^;�cd����'��%�<�k��q���$���F-1�;��m3�'z���aդ3e�F��tx}P�ݝ�.�Ӗ��DC>k�S�̓�L�4�s�L��t����,�����׷6"iPg���8���$����NM��HQKָx,勨>e��=�d̻ۘ-֛;�<(�Q��_����U�8��#6ƕ�]��kf�ri�CqEc�Y����И�/�M{Z�E�&�{�l�B*��1�����L=�U��.8z��E��2vX8n���4`yiC|�h̆7U�'QN��r,����p�".k5�5n���ܧ��R�S8&������d� �M���,��ob�v��i�y��ܐ������E���+�q�S��\�[�d�S�&�7�����Y4�9�R�\��4FD�pD)m���҃�xE�Z<}ט������k���K�%f\�/��ʩf%���R�D:�5��HЭ�t��A�*���;ȳE�5[�������YOZ�L��
��t�<m�� ]���K'�ߊ��w0�3C$�cn��UV*i�0��t�z�'W��B�Z5�|�=Sp�Z�L
�����{'����ޟ
L��\؍9J$���?�p}y����M|�}~O-t*�W=\V��:��h#5���T��k�=���HR-��8���5�t��Y�X�m�	z*��w��P	� }X�XF�f3T�m�.� #�E�#|I�˯�k$�\3F���R:4�z�)�%v��έmڙG��5S־���Uj�Q��Ki��趃[OϿZ����^tΩ@��/Gf��D6���7@�S���g]�����Ulw]HOlZg��L�؁�S�LuR�=�P"���y�UE��H��Ii��,�-� $q�A<`�0\�u'�AȘ8�4]�7��z;�A{�X���򹇛�j�s��<8�R����Gtr��q��wms7{ܑ�26��kn�bѣ�S��9��*���%ݑU�D9�݂�)�Y^~a"EU"�)����7�
մ٥ǳ�d���O���x�a�qW�~?�B���u'���G6.�����/�R���D��	�㸵^ίf�1�X���%j�Z�:��%��� '�\:C�me��*�D	�����ۄ��v�i��U�G��tS��s\��ߴx]|���Oh��c�pU<Z�G"?l|>���UN�
96��^!R�qJ�7���S'i���.g�|�Qa��!�o�g�	�ƕ-@<e�Nho����`��M��Fa>��ϼ����CU�M�t����k��(,�8�Z��(�%C��g�PO$tF�i�����(����
j�ǨW�7MU`ƶN3N-��u�I��g{L���Y���c
���>�Ũ/$	/�>�𳔂iE�y6u�RMu�(����M�Yن��~�]3СL�τ}�p%;S���ߏ�o��u��~(�hn�� �X�Λ|,�>�Hрu��qԴ%<
�|e���׾fn2"?yz�HA�#b�"��ŝ��b������Y��Q�~O_��\��11���뮤��N	�rz�־E:���6�>�E;�����ـRҊ���ֺ�|~ha�����W��<q�,�Ȝ���o�P�⫔�_���G�-N�a	=�Q�Q�f�l���O��X޾5�Qˑ���Ԍ����dn����&����R�-y�?���S�3���Z?�#��xZK�O�Gd����fQ+�Jt�����풠�S.s�Z����?��
u��a2đ(�����7P���fnbq/}��L��~��sʳB����tjj#mSX	����B]�	���n>� �d]p�~�2����~1)ֱ�k_��=�}k:3֤�͓_�_�����fP�t�_���5/f�h��xe,be3�HL�����QWb��l8E��=`����x��a�^���%Q�U�%���jzw�'�d�PG
��B�����yZ<���|*	�ˍ��q4$����ֲ �� 10\�|"����1����B��A��$�9c�G>%Ee��S6��q������:�vh���V�C��WJN�+x3S��G��B�߼j���g��~ӓ��Kw���y;�>~�|�����2"7����F�^A��ɜ/k��u�:�L5���=e_D�������:g6�*���� (~��� %]�4�Θ�l��u����H�S����`C��0 ��I9�#��N�$'����mkk@��;hH�O��q����X� ��([^(!�}#��A�T�y��[b�~x+b������AJe&,A�A~:��������g^r�1�$��i�R�Z6�i��%Zzn����G%߀�M���!x�Lη��7
!�׵ᚮh�Z��)���)����*&�f|��ɾ���{�l�]��a�u�������([8�P��j��R1��V��%�)G��H�~�:��՞$�qtE&c��{�0�Ь,�"�O�;�����쪪1!�-�����xIh֗����{�9 ۪�=9
�n��5V�By�&���f�&��l�aAM'ӯ����۔�^s�����k���g�o��|��BaWP�[`l�d;l������"���2�G>c�Ls���1l�ڿ�{˥"��X��"��ΜJk�([ B y��Ы��Qn��΅���2M�N���f�=�Ya�{"%��Zd�
��'�׽�8JPc2n��E�^ڱM�
��:�gǵY�ܵ���TĲ�F�w��2PD�+���Q|��q4�c��2��,n�}�r�4����$s"		���A�����o�?�j�E�k�����M00���:��8�wݾJ��ih����{�h�˝н6���1i�D�.�'�ǽ^"_;�
�O ����а�����Ot?�^pwV����\���n�?��,���A�t^��G榻�u��j,��Oݙxwsi~���P��GV�����]G��<NX�45G;������Eʒ�hEVWb�B���Rӝ��݌�նZ�]3Z�%&��%��^���?�RY�����}��oeF��)A �pa�KA��8�L����p�'��6��q���ρK�O�p�sM�rP^���䋭Ƹ�� ]�rʃ�5��|� !��-$����5�L����P�c\Y�*�הZ�!7������f�j~��^d)�%�?�]m3��u��`��G���pv��|�Z�c�:����ۙw��t<���E�ɩג�N��z���qڄ`� oU��ֲ�Դ����{K�-�n���A�;H�"{pC�ma�A9,G	�J���kZ�ӟ�x��2l�5a�F"ċP��~¥�
`Ņ��|3율�I8>w���8��������p3_�Ց��)��{�
��{�h���/���������~�z�����U�[�G(�,ɕ,��Ch�GyQ�|�k6��f�}��j�?I��Q>����#�t!y��%��7��JƁ~�R�?9%�D�
��G�pUev,�T���;,Et"@ �ʨq��Z���Жu�S)~_���A�e��m֘k�A���d�J�$�湮��#���6��"���a�|~FU�[�#{0�=c�;5`�V̝�����Z��,VC��{V� ��Nז7�b�V10C�Hc�0q'�&aD�{O@���o1yA�tN�vg�:�|8��뭩�8`��n��[�d�~5ޜ�y�_�v�32�K��u�F�]�s�rH>+!pY�}���������0.k�K��4Gy�,��m�p$�(���<�Vm�|�GڼKX�X��S0���QR�Q�ӣ�u�+�0�{�ݩV����Ē�{��~~�7w�Yj�u��p�UAǵ`/��@P{p�;��TDx��ঊ�'���T �؞�1+��q�����;���O�cc�<��eg=i�^��۩�����_��j���I�tJC��D�㼹���I;p�H�ABOa����d�<���������̿y��\��U�i�sޖԺ<�_@,�L���ͣ�p�����w�]S��1� ���f���_��Nˣ�15����5����>0�0�^~`�-IK5���,� N��Vu&}� �c�+����l1�i�8!,jwY�ɜ�.x��̰K�\����ȣ%2��qS��a"'��WM% �P�F�?������9�yAp�,�
B�`|x��S�[��D�X��ӧ��eQ��Q!�Y��.��`S�e��5S��� _����9+��d�6])q'Cº&[XiW5�|�Q�=�*^%F��*	k��h_#v��>*e�'Q��(dι��]i��/�yl�Dr��˛�U�k���+��
���>�̺|�;Z�� aӖ�#C�,���s3!����4����-x�X�y�Ү����D[��}���y�"B��XM�nf��7H4�K[��\Liqki�̒r�y�;��OHZ����,����ֻ�a��0o���aZ�G��[n���u�}o5�~W�v})`�СХB�>4LS�g��"%��$Ul8�U��M괿XW�x�1��w�����?�$��'���t����������`jP�w��9�k��ܱV�>�2��lo�[�9C��C'U����UD|+�;4-��\p��%6����3Z�;��l��p�p8ͿZ���>+�7�	�g��(����c�MJ?����o��XvϟJ$�Z�`��z��<Ax�<O*D�vx�U�{B�UV�p�^��l����O�"�f��?��u��D�V����of�o��k�����B/����'n�Q��Ӧ��\����2����<�r�Vs�8�H���&C��ݺnʔo��6т��d
��|X�ƺ�|�����ce�(n�ң��\O!RLmʙME��\8y减�1��`L��)����t�Z�EUɞ;��r��g���Tv��½d��.b�=�����"8g>�ao���u ZT���dr�iL_�\�r�Őψu�v���O����޵��/nIG �'�����mv�_H=����ἡy�Ԧ��	���k��Ӂ�Ilhd���{�n�`�H(��d^�@��5# �*�~�pCD~�LRr���ɱD�\`^���v ��]�Q@��~n �o[���n��oH��_f���J>W #�:�h���ʲ�/c�X�;K�z�|cA�R�p���q�4��ʽn���tp�v��N���7�_���(��Zm�lQ�&f�\#� ��P� >D��B�j6��%�`b�=�< �#��Ũ�� ���|�t��[��C��y�	�F{3�M��nj�O�U-Dy��?�<�~.���r����5�vH{���>�p�pcFa&w\RQ|�����/͟2��"�ZDL�����Gk���6?"���p�v�V=��5\	%3D킀o o�>�Z�YP��kc�d�E�����©C�C���N�{[*�0�f�O��L��>D��&p��jY��*Nl��/�'����~
�i��+BIξC�l<�BUMG�g���z��#���*��o}�/T�ٻG|?�7�r����8�ݦ���@zM\f�h7po��3
� #�%
�v�O���2{]�,ש��=	"��Cf��<�P\��ap�%���&���㱢.̭8���Z�F��^��k��Q�FX{�����C'Q�]7I%lK� �9x�l��P����4:�s�Je8F����R>U�F�3[��1�F���x4#I*3��a�}��Z��";�Nn�#f������DX����ɋ��s��Ro�z��1�݁�4)(�}����̻F�S
�ȗ�rJ΃�%�@u�m˨�E"PV�W���~Y~�5&����N|��������'c���E0����l�I�C�;C�l�-����*z����:Z�7�^=L�f��p!V�L(��8�����XV�ci�_�Ɛ[7_Z�F� "���k�e#%8��1[#9ȗ�ذ�_��U-��Σ��@4_bt��}�זߎi�@ f�[N�!�>z���Q�XYd��z�G�Em�jV��=?SZ?��&��N����~�
*ɶ<o��̛�"ݨzj�g�F���Y#Ԇy� Y��Àd�/�i���8�yh
�	��~�ꐜ�?���I�o��W�]�"[c�yA��p(��\��ޘ<����A�:�����m� ��I����J�`j�Ɔ>G�B�.����P�Ċ5�}N��Uil�*�o'���3�#�ڪ�֘Dp	���:2�M���(�6e�1]��w�������GZ{?1�+��6�ʁ��3�Blu�	q��Ҍ$�,�0�8 N	�� 5��oG���a�����.������	,��*�g�T�����]	�k��b�Ts2?�߂f��k��yR)]!s���S5$9�J��%�F,�ҡC����3��]N˞��@@ ��7�ap��<�N�����Дwx�@c�I-	���}5Ʀwr9����乶�pvYC�EÆ�)�I�vE�.h��������Ɉ�6I�{��WzN�N}�d�)Cv|5�S{�а
����i��(rϏ�n`n�]=���yc�MJO������$��e��?5٭�Sv�
'z���gb�2yiM)�~��W갖9U�n�AC%����<$�Έ$�G6�s��~Iy��.0w�>����+'^Y{�F
��!z�}��LHU� ��K��#��xP��T%�D5��iΈd�:r�hJ�62�{��]�1������&��1�HA���y	�p�e^�D���RQ��,� ��W�Shw[`iܦ[���M��!�����K|��Pҳ�)���Y&�:�D��������1<�O3�@|��?6��!mK4���Y(|��(�t_Z�|n�8P�r�#���c�z��=���h�`�zPQ+����rʙ������:ewؗ�=�ɿ\�ch4WB,{������MD��� �|�^����E��R�cI��cݒ�G������'��]0H� �
�	�B�Y�ej��XZ�HVrY�����umv�.�᭾1H�ޤk���y�M^��'�8��NfQTS�h�ҙo�8���*�F+r37�jղ�5gA%]�!�N��N��φ��;�7J!{( ����ͼ�-�(1g�����\����G���3��O!���G�U�Ѷ��>�j{ǿW��L�����UG��z��T�\�����vlIwu*6�Q[�{��ܗ�Q˲>NC[cH�q|BsÜa �@X<6��Q~(זG��JW���C<�ú��~�~�S^q\=lW;�r�8o�"^f*�~�j�״z��2�(C�w[�`2��=G�cl�O=���)k��43$~�8�P?��&@GZ��N� I��v�eH��y-0�0Y�[�ݸe���h���Y�"��V̥{ׄcq��� ME&�H_��`l�[ڥ�=Ü'���Oڪ<-T_�����} �A$��C3�z=��9[������6D
(=��n��~"b�c)��V�^�������kB�GB���r�:x��uS��&fn�!�͟\��97f0jP���!�aF��r�0 k"H�6�!�����z�~���I�N�Jz��%5K�%T�����GdԀ`�!�-����̀���eo�w�x*��k�V�����v���8,��ڈ�kFy��3�H��RWƁ�[ �4�ਝl+u���Vq~���j^h;t>Q���m1�a�v�-/�1�� 0d�����"��o��0�r��m7q����s8�5����ܧ[Do��Xt��p` 3��i�؟Bi}E�x�@|Af<���W#_)W��S�����8�`{J�|��ٵ��F ɽ5`fw;����P�Υj�t�?��G������������۩B=�+7Q�E���d�Tbf�Ѭ�I;pfN��|��$em��P����;��wH�:p��8�QZ���"��jp��'�d]wD*���=o��B̔f�
�I5'	ܓ��2A�8�����* ��PǖD��h��+�-Am�D��H��x;A#`ΙQ �������1��.;hj��F���Cr_���0��|H�e���(�R�0Gme��cKW���q�Gu]�T�;�}�N"�FQ�)Y�W�v7�l5A6����Ļ�yvʐ|�h5�i�|��GI0^����-HR�NMM��O8� �7 N�\仴Í2���ȧ�/����ˡb��q�z��	�L����ߨ�����_�g6^U6����a�u�U#���-�T�%-dp-�P���M�9S�=����ѶO.HR6�O�eJ|�w��8z�f���4Mц�k� s��Yƹ*�б���&T�F�y�Ig+E��:����|	AN:�}S�S>W����t!�N	4�v	�P�ͦ���O6�]�ҩ�!�aڷ�|W�y�t���d�f��0���\0�b��(�1�it�B&h6.Ƚ؈�
>���wC���Q࣬�*\�YSG�����-"R|��e�B\�͖��x�j}"�`������Rq*7�>(��w��S	��7��pe���b�x?�?&�?g����$Ǜa��	����u3.��jpو��O�Ȃ�������vZ�®�z]�w���;>�`f*�����f(��ѷd/���/�H��M�Ե�	�o|��Mo��X�[ѕ�',������ &�D�u�,�q�J֊<Dgb�H�dN��B���=����+%=�}|��$���_kg�m��_�-�o3�Az9�i���>�!���F�@绦��4�j�?&���|��P�X+��Ȟ�M���aC�1���{7* �F�rp�O�P�����ab���>d
�{�=[퍳R ���%�佭��2�����آ\�uaV��Q��F<���
��'%᱃�ſr�	^/
.���W)����2���4k���X����pm ����t�Ohbu;��\��<�~�?ג��Y�KH�d��"E��E4����$Rc��95�ʲ��]��Ϊ��+Q2�i�.����&)[s�� ��)&Bu��i"M\7 ���v̨�<�T|F��R���"h4U��b�'�5��ђU��nZhG�F԰ӑ�cWyO�&ٿ��)h@�`�|
2�|3��:f��c=�;��@~̟�����i����٢/��ܿ,�v蕑��}!�DUV>��/�C(�H��E�ٟ�`��)+�!K;��'C�EH�;��v��6��s��l�w��
4�Wvc��=�y�^SNF�?��rgV=񚔥���s�90���#�MT��3Mǰ|4�8���t��˞h,ϐ/�/�T];+F�K��(X��H�fw��2d�jM��Ő�a��H{��F���/�f�'N��U{͗Iϯ�U�6��\�N���s��}��	��yw*��b��H��������9}����Cn����#�u4#"ܵd`3�^��Ҭ��n	���,N��?��jՠ���5>�|���D�C�zū�`]��C�2$����U!v�!-O�z|�c6�f��k��Z���$ �,���"\�����De���.´{�����j3O�k� ���5�Z�_����Y�9�տ�` ���Ȓ��ilQ���EA�e7i�����;<�<볶�;������wU�81f� 5Ns��r�5�S�w��<��:+]:��L�ap�r���w�W\B?�%�?Բ	��&�!�@�Y���s�s�1'�iJ��B���Àq��X��M,��<����P�^���4?����L(�p�r -��]����5�<�U�;̢͟0���� �
;1���_�fe��u�q'q�0[p��|M{j�U�\ׁ���#����Q�j$(]�[̽��2�V~�'{��i~������i;�LQP(_7$s�N��Q�8��J�\긆`C��
dv��0m6�,�J�9��ה1�K(�c;�^���p�kz�?���.a�q�]-�����G�f��C�︦�@m`m�rϪBs��Q7Tk��=c)m$^sx����ʔ��egMU�JE�(N��E �a+fL�T+�SʣЗ���t���d��/p��$@���=&<_��R������$��9�~�|8U������Mrn����U�"m�Z����C�xs�������e���LX�Z�1�����}!��Yf��p�󏲴��� �P��9_�c���0ա$0�r	s!��4�kh�����m��<	� q�Ճ:+Wp�XRg��ɃPX��?�\H���6���q1�����]\�k��9�x���Ҧ3�bf��-^T�a���଴��	��D���V�_*SC=����2
��g� ��N���\�E�DX|������㴼�v
p�T~���M̦,bY�1�¶�\�F�B�!�>,�5(��� Up�̼�3;��ކ��{͒A��g�ˍ�BR�p$4ݐyG�kL� �R��o})}�A�k�U�������_4є�C!�
�4aW�F8��4�^~��]M��3�_����b�ў�Aϊŋ��v&�UAf��.o�1�bo���3*l���,��g�ӿ�FP<$�)��w#;���貳;�x�o1� J�2n֌{$	�%��&.�
;!e���P�%�����D�����a\*urx�'z�§���5��d�j���'�	��8�(t��Q�E��k����Nr��z:�������NQ�w�u��B��,�XY@-W ��\�ם��`̉������N/Dz��/UMˬ�K'�&���xo@|�]%�lr����J�P��נ�5O_ha��������Z����m��zSH��? ���ɌJ$��[K��s:`��-S�b%Fx���q:� z�������A�B�w���I}ef÷+;�\�͠R1��)�c�+�s�X��6EBc���s�T��J�MY�(��H��iٌeg��fb��$��|!��V�,N�����Q[������y�Xm
�N���xvs0���Z�1���T�:���d�M��-�8��?o۵+�hiwŲ�n#�e1m��
�Sל��J��v���ў#i:v�J�~,�5��{��ࣤ/ �H�ۮF�m.~�k¼�>)�=q�h\���nÒ���� ��(�YɌ�e���Vy+-�6�AtM�R�����B���/a\X����]���v?�,p.�����T�E.=���"x���<�6�(����p�h?�V�_p���1a����rї��g�z�qj(�;p�W�)����\T�%:p�0S}�b���"`��.?�����5�i�m���Y�T�q�g�����j��:�y��f�e��I�SP�[16��ZK~凶��P%��eo����ө.�N�Z�+V���_�`��։-�Z�#�ς���.)�Mo1M��;]����웓��	F��y3;��#������%���*����D�����l=k�t<*
��Ew������p ޶3�[��t�m'aa`�RV�y�)��#q�K`��g>Zl���͹#?)Q��@�)����IF�]�Y0ѣ3�QE ��p/r�)s��3J��W�7`B�ߕ=�wfkqǹ�Bz�F�e2�&&Ѕ���w�eQ%��K!e����/|�Y�5�|DLÝ������̸+3g�2y�`/������fͰUc�k~��ꢎ�f,�Ҍ
6�&����5�㞐��O㻄�D$�z���=sF���C\��z�v��G��z)�l��io��:�ޠ�`Cm��{��a���Zg݉��n�;X�r]�H'��_�Z�f�� [�S��Bz&�؆��=��$�X/->��� ��$��('�~�<��no��h�+MdD�,�iS��B;�Q�"�_�o(%G�넱������Woa�z����&�>��X��:�f؉�7�|0����qO滕Cw��9P7 rc�2����߉\%�;#����ga=d���ۡ�W�z��,纨Y��6�!�?:�e�l2���hA&8/��>j+y�#	��2Gtr{3'^�=J��5����rP�tT|+5Ir}�� {H�?�Z�jc���E������u��o�l���_�m9Tٜ�A���S�r;���[�Z��~�<*�i;����0>�wA�S\�W�ZSΕ*2e%>K@�.h�eP�v�Mj�@e���E�����ѳ�FV^�V�>�1� 'Q��o@�U�Px����	d���	�A����9C����[+�j�%����o�2�d��8����~kb��W@��h�u!�}/Ԓo�����zU�.��l�^\�\t��VN}i�6�����յ��!�#?�Άb��� ��C�08,��n/��V>-�@Hݖ�5�,Е�'�E.G&:'�"�3�U�_d�?���M����㊷���YEm�0%�v�lx:�]!���)�0�Q�����J�'r�y�y�_'�]R)nElzfÚF�a���	q#�c��X;�3:��֬z}}S, ��/��R�?��������x;4��1���R��
�1�-=��&���>$uGG�-`���=�l
�ٚ���
��
%a3e����� �J�I���rnsC���#��v_uBQ^ ���`<�[T�����oP|c!t@����*�������|r�2�X���"��%�:Y-���x�*,ϱP�w��Gbԛ���m���#�KuE�������<�U�~w�)}g�y.�Ϳ����R�!�I������)�f����i־�t�#��!��e�ѱM-`�vi[��f<`V/�KE0�Л�B�2$�X䎄P�H�]�~��^���q����Uȁr�(� �lG�T?��≠��KdX�����ؚzDq0�	�T&eq?�,�L�ɮ���mA�è����oU��>��JR�M����0J��F��t�M�^>̢��hQop�لV6�P����M؎����
J��.����O��[�?�򠆖�he��*n�����{HZ�d=�p��B��`���um[~IS4s"��,�0��R8.�i)A�3ӈ�K��[&BP����&mո�2�X�B�c�`���:s�m���œTN�R�%6���(_\��j�3�ک_uN�B1�[�͠��p�ҤR�����(Cz���)�+��$~�5���,�$��)�f�\�����e���0�*ƹ��怈�%���?�Q]��=e���2�8��]�6��D�[#��qc�8��MwS��_c�����ɚM�װ�������$�p!�ۮ�v�3����|-"ɽ��z��PA��6�jGf�wtQ�G��M�5\��*%��m����zc$���:�!J�"j� 
D4"�����#Ǻ��r��neC.W�/�IԄ��mM��j��w��ݧ#i��O���&E����������
j�I�I��fh %�ZA37��z���lI�/1L�[H�#�����*+ �<������D��ρ6�␺���0�ZҶt�RXɸ}�x� ^�v�V3��,ҮB��&A}�R��ҧ��;���8+����8ӸA�&�x��$�.�HIT�	�=�M�P[
�r%�����r{=��%6�2�=�`~㍟�'�>�pe�0�sd޶.�H��`�����ͫ�2=�T:���8���XYp�wWt/�yx�{���	�'h�ʾ{���f��1��4A�҇��	S��1y�^!�v�J�@�Q]]��3H^������!�Kr�w�iޘ�ϯG]ͷq0���A���8����#'1�Լ|΄�u��������ƹ1g]����<�Ԁ��2{�I	���U�zKo��^VE�	9�N��:5l��1s�39�M���e�:�X�z8@�q��*���A�W���:��e���\[B�U�����O��"-��0B�)0$+�m��	��ܔ{C;��CZ'9-��3/��C�28��hA���q5�`6���5����i�Xq���)C͠��:~�[Xy�F�ҏtV5��w�ڪݑ���>k}�O;�Y�­R��<k�F����7J�#�� y/e��;�[��8�A��@(�`y�o�	Dc������֖~�� ��ƶ�٩�x�@�P���#�M�����[r}��P����:��8���g�8�x3�!���z)�-��+ q��r	3Q�S�������՘����D�pkå\rrr�!��q�ߝ]\�^�(T0��0��땡�z��Y�*9��=���<'�0.��b|Y��/�A�	��9[�͡��� �/͚�;����_�������yw����3K��H+��AZ��`�8I~��(Wi)!m!�������Ab��Q<�.j��أ�}�?}��*�Kz�:����l�l㨓�̚���F�6��C{� �3����џ�`n����v].�a��������k_5OT�e_�K�?A���P��+�\$~B�����?'������p�%��������aA��ے��>�F$�	LI�Ko�+��u����8=�*�땸�<\�%��)N?�`{�����;�-A�@�:�� ��? �^%{���C���J�c`3ݹ~��t�H@�̨�wC��A�d�ʎ��7敒擎~*��5����8�eX�o}m�.�ºĢ���C���=<+[������2D�����L(L>����)q�!��<����U��F�(jM�/ >�[��v��XU��>B����M
�p��}�n���Z��F���{V��)$H�hTJ���vĶ"Ѐ�-/P�23�Lm�^��E���a�J���O�! �'���^Gp�1�a6Z8k��?�
Λ�{��F��@P�l`2nkmՍ% g�0}9�؍U�pQ��t��[���q�@;�Vv����I>�E�W������ҍ��e��J����2B��5�4R��V��^6E�Yo�Cn��=�LJ3���S��B�B�yBb����@dߍ�ݘS��etp���Ʊoyh����K���H���%I��_�6e�:�{zCUY����H��G�4s��F-Ů4�q���%�6�Ѽ���|s%f�ǝ��"ϑO�e%���3RT(������%��r��B,��jH�7d��U]X)f�p�$л!�S�m��3{�X^�2e�X�ypt(��"�Fl���Nc�-!(z5Y+Q�'��\Vw�7�>���"��<#]���X��X��g[����7��?�?E'��q��I6r�}��_w��������	��~x�o6����BX��L�{a��G��7yZZ����o�N�6,�Z�F�}�f|��8s� {�N�� h�j�'��<��8A=&�x��M\k`7�6�S���9gnͽɋn���HC�Ugf����1�B��J�]1dhF��~Ʉ�\�P�N]���:����EW��(�����įt�^�s�>IrP�0��Q�wkp�M��<���P�nmn`V�6��ӎG���K����p�魷k	��k�Yf�$������������e\��iQ�S@��Pi��V���`.>%��6�'3����;{F����1��d��Z�.GMr�86��2���ݴu�ژ��2R�"�����d|��U<|# rT��p�=0� �Խ�[0���͢]
���R�rdd�7~xX��1���Qq?V�|�=R����k���r	�������2c�$f$�qm3��ԓ�	X.�Sg]��(ߓ3zg��Tl�L��$�XtC+��D��~�0�A�o����l3~�G��|�6��>QX����Ie��3i��(�>!7��Z�ku"������e�͑�1�:��v�n�^3.���������8B"�*����r7��΢U����_G�2�
cyL�6V�)W�ƊZG���T��񂃻B��
R-4I��AA|C���lՕ!G��B����5�u��S���g��>���8�3orr#���������r���|q�>L��wmm��:��^�w	D j�*Sč��P̻�3�/�)J���J�H�R%�u�/m��O��^x(cimø�,�<���8S�ۡQH������<�1n���*ʓұ��e�l: �R�8�(K�pm4펫��`�ɻ���Z�=�O\m��|��i��i�X2:��Mp'(PV��ۺ�7��V�U5h�n�$�Gq�s���ǜ�ڊR>���5��������v��Ν&�iZ��[%��%�I�:��@�=<��J����	��g��2}���&m��3噞��kӯ��؛�eV���#˄��Z�fN���̇�CL����5���1zp��7D�d]؃? ���Л

�3І�a����}D�@�J�@�ߝgd6+�0�d0;�2Y�=��R�`v�|��y��_�T"1n�����*
نgUo���"�.�(��:
��ؖB���\��?�-4��ވP�u���~f�^	�˪��2���l6��	�������΀إ.�j�VN� ֮�;���5X�u(+���RrK�E�_L��
�I`���
<�I$f���Z{U��F}VZ\�@^S�>
e+~g�(��ь�J�\o(��C`������6'��L��; ]O��ԗ6/7��6q�ܥ�뎟��x#LHT�õfԻ����:(��
xߔ�X
}��N[�O�ڦ����+�����?�?T��4��#j�I��Hֺ~��>]_"������\�\l�$��&E;d�%T�u���p�\��K�A���|��.��/s���KB��9Z�3g7AX�/�5S��}!�����6�^O��jܱ��G%1�z��p�l~i��3ͬBu�p�c�.��Ҡ[a^�s�S���x�9L-�!��鳗�5����uV a@��N�sqtYnm��u9�Q��ԭ�1-�|R@�l����G���O�_�2M�H��q��emG��ƒ���j�/Aj"�5,>�,���:��D�z���a��Z�i�
R����7�P��D%)��4U�%Eʇ	�����^d������dbs�T��;����ߦ�St��+f�Ƶl��Z�?q9̹�=嬿ݿ����v��#0V��{����� �P ]�%�N'j�(e���P���&�d��gFD^F�Jc�ǣ$�`~�<��Dc���9�\��kqP
��ao��z��X����x ����)�jZտ\��ױ���b�[������N
�,�W(,���5�F@x{�B-�
�6F�)��,�� 6�$�Cf>=;�~�%�u8*��ǩ�?v�_�ޖ�* ����'�-z��_�P?�1W�3M�k��(�Z(���4:�_�Rw�c��}���3���S?�U��V�$x|�	�J�זC��K�a�?�j��z���6U�=�nR!�yx:��c|"�âF��cr8%n��'�,ꝶ'`\M4��C|�87�Ǭ�����:ًWU@�����A;�\�7�7^>����O2�Y1^��y�gn�ZT�/��Q ��
���� ��R+�g{j[�#4͕��݊#hK�#�HK�9����|-�(����R�ϋ t[gd���Vf����-����h��7^�Ac�����4�@ ����xd$��53���F��w�!�@��H@��|��e;���Y������M��!B��?ԣoҠ�m�����lh���h=���wa	?k��Yq�<h��F�^��E (|;���.Y��N�����Ad��K��\��QPT�b��s������7N7�H{���׫K���ņ���$Xj��G
s�sWRa{| ��y����Y��Ӆ�$JXn�r�n�+��'2��{.D9��`�[#�>���:R��'޹h�/��m��hF��G�Wq����Ԇ�,C{ό��&r^to+sBP��u�b�����5Ǟ�&��zf����hWPzˏ����S-�|��o�Ѐ��)[e��bTdKN����
)�����ho�w��D����E�?e*�G}�mP��	���N��}��نn���e˥y�O�1ɢ��򛈘E�_έNv�p�f�a"TÒ6��8aƱ�Qيb�2⽽?/4��|�%��������K�W��|-}�>zF��g�~?G:%�7�BYR�c�1 �Z%����d��x��=:]L$@�ʏ6N ��1Q��=��ب	�3��+���ST�j"�}_|�����5R�J��,�Bc���p0��Ӓ��oD
4p��v��u��?�BJ�a�#��M�耏=�c��u�`��3�Y�Q1H���/����ܵ����:�7c �jaJw�`� t�� �j�C�Ah28��^�\�40�Ԃq��1�6?��<s�j�-IB\�����$���۲e����
��G�� k\1��[gX�Y��W�{�ٕ�{F��1���������.p����_�?��q|[����͔�!�� ���#�'����;ڠ�����%�qH�_�ǚ{���k�x�����b�:�pg��{������T�{Ϫ9a���0A�n�0�ߏ��
z�\PM_�ܖ�H.�YK?����/n` k>-S����L/�> ���G�'f&�=R�Z�'�Lp�}�#bo�����|o=(�=�~z�dqƶ#�k`���[�oG�ˏ��ط$�֊QBF�p���OW��Wb〟�f���#�|o��G�k���l1�4rOi�C�-;Y�[������|u��G>�H�;ŭw�j�J^t�4�m%�{ؐ���[Bp#�*�_����x��j�}.+L�,{ϫap�K�˹W���wn� �Ѽ	��c�H8��a"DM_˯���3�3�s���2:)5Ĝ�Ɲ�x�	o� މ�8�wP�a.~be�.9$�}���+ͷ|�^ȿR8��ô�δ�e���P�f��M��"H����/l�1�&�*��2꣙�`q���S�X�WE���.F ��S��H�QA�^T�}�`�Ț��匐�P��u�?����2�<��qOY�X�D��dzɑ@�oU"�ވ�Uj67:"@��βQ���6*��`��@��ͽ����](2}�Z\1܅�*p�q�oY���|����+E���3���rag�]�#6L,J���r�����}WzT�M���K���=����6�2~Op�FX�m��-8LA�|Z���;��&IO)� ��j�c�p��#m}�}!�3�m4*�
�Y�h?푯��~V5��8�=�ܶ}�D6i4�� ݙ���Ot�ΉPv@�^�oY�!�>"c��P�Ƈ�Qҽ��7�������o�	�@!�K"q�@u"�s��om�Fr�D��  �@��cUKN0��/cG��;P�jx�PKo��������,�q�vf�N��r}������s�HU�1�@���b\�,���F)WGR��3����j��+��ˀ���0�u�H����V�͋L�x{��Y���`l2ʊvۂL���]s�T�C�����RN-
�yŖ�܂Ы)�%3#��*��m@Н����b��}t��9p���>=������_�t.# >��x@�]}��g����

yB�z�*���t�/�$A[���
��1�DHf;��cy�P����X��H�/�ዦ"5�~��<�y�h�wϴM��c?��*+T�)E��Z�gL��$�d�LM�k����Ǟ�Dp1�ֱ�k��`��[�Ž��;��S��������g#�������2=n[�{�{,2Q���{$����n�ݵ��΢�������q�|VW�5	wK��_g���L��B�K��I1㨤��d��YT�껟���$6�0��]n�6 �0X+`�y%*�OAY#�H�!�F��ĭ��\ca��*�E���Q?�C	�a��e3�,�L(	�US�jq��A�)���d!��t1��\��1|����bI����lF"�꬜�}4&������q��R�?.��9�:\N&e���o3�P�J�)w��r���`A��p�j0��̳��M��Ԫn����yXDtᝥM@v�7+sa�̊���_�4�N��r|��=�.K?s8N�y��`rvM9J51|X"��1��7O��~�<hB�w�5�j��|��
�4�U.֖�JB��1[~��������2�ބ�XF���E����F��d!�e,!����cl��ywͣ���� �l�L0kN="�F��4��֏�-~�W�'w'py�����+����⇉���׵u��)E�(1�A�>�q)�A���n9vD�P+�g���b�%a�\�b��RN��S��������r�l�)W���P��@�I��A�Ҩ�?�����c���Ԙ�l�D�.�̋2���:��x���&d���i�<z<B���b�o�<�)ڻ2�L, r6�6�Q��R^N?�5A�>��~x�ȧ����h���-�ԁ���ߧ3���Hr�9fY�+r���U�w�o8 ��@�O�'dn�s1���%�=�
�;���\�w:r俙�0vb7E�c���DZ�P5~sp���T}��;��Wt�>�5PNIJR;-����jy�����z �6�Ʃ�!�#9p<�?��%����œ��?��-@}���d���Qu�[�T)�+�̾�F���'(���
e�x�p�BDD�$��*�A����
��g �����@,��3DN�;��B�S�H�^+g��5Z.�|�����[p��t@n�:&rMD20����ᚵGZi���W���ʺ�wY��w�uy�ň�im�󸩿l~�G�`GoMBH�:��=��YL���[���`���:��5 :D�̃r��LM���O���?C�3�!��4G�	�Z[d�wTR9ⷚ���1��=
#�cG�~� ���j�G��Ǯ�����f2�^����}2�έ�> (���z�K*����;Ia���_S��O��J��"�&��X�z.'����Gc���;�i,����mxW������ַ�MMs��.wNF�J�l}:Q�2#N�;�рY|�&��@/��3*o��lo05z��2u��Fz�⩫BO����M���?c.��Ɛ�<QRJ�x�i����� x�ǹ��'<Sӕ_�e�Ͱ��˶'�=7N��贈^���:�O��O�'��_�|Уh�#FT1�uL-�<�)]hq�UB����!TցSx.��	a� ��DW��;��Lkx����`-\���?}��IP>	�.Th0��.'h���� TВ�*�|��e�	�@�p�̠jK� �9
�=X�h�#K���:I�DF3{��0���|�Qm�絛��5����.�St=�`������+�,��m�B�)�'�D��S5r�wP�<���@���+��9i��W�{Gk?��;�|,�4����.n�93��1�~�m�o+�_�&�K"� �vK�8�p�����X���<�1MD��[�+�~�Mc��/���M�+;��ƓI���/�r�^*�Id�-�7�u�]D
�׾��}7�~�[�j�����դ�B��T���9�#��85���.\���:l��n�:�šmy~%T��z.��)!K���OP^� �T|�4����4V:�͊��$#��|�BP뉊�a`؈N6u�V٢I�����*����T`���2���\	޵؋�}��.�I7���L�E�<����3��>=�v�s��\6�L��QB�Jcf%��>��@��%�v���1�z�Y�ä����\|�2�E��W��H\t���n��cg#1���ZW�[ ً�'b��6FZ���X7ћ��cuX'���ٵ��B�
�a?omn�f�sk�t��߳�v2����ʀB��i�Y�;ʳ<B�W�TP��N+1Q�+uد��y�t@��������$z�=�ژ�nx����&�M��~C��e��dgvC�y.>���.4��M�ۑY����u�?���A��27E�� �� �e�%Ej~,E+3]D�О�@�a����<�D5��/�ǘ@��i����{��F#	T���,��1^̴�zTD�(�)k��!����hie-�?�ވ��~�`P���V�kd�3�p��
��Iʪ�&7OГ�C���'6o�ǜ���x�=�ct�#�t���7�.���Q��ᡯwu����@�$r��P�t���:���['���]��_���mDfo_"Wgi9�0�����i?�#����X,�Ŋ�$T�N���?������R��2{�xfm�ᰠj¯���+]NJ/�K%2FŢi�U��qԹ�Y�>jFa-GD'2�*�|�����J��m���S��;�*�|M� �hS:�$�>�b"�|�F�w��m!*G��������6߯� 4�H�ڰ|�܋ۤG+��Ȋh��۟l@���5��N<iuAo<	�`��6Ix�OHC@��l:rȕК�y^:� �{�9���/�f�He�Ӗ��Ǳ/qmZB�����{�Yp����~h�:[�Cd^?��d���A�v��P �
�ڂd��P����_�Xd�.��(�5S���s>�b+�b8<��e�>�B�«��2���?��Z��C4 >c��y�UU��B��"t��xȢ-���G�@7�i��C�쎆�q�����-�����Ϻ.�Q͠�ԧ�;���\�m�fU��/@DG��wܶB>*5n>H�t�K��Xwߟ��R���}�-׮�3O��*�k����̽I*p��]F��+>:�d>K�#��"�G�+��1��%��ܧ�WC��׍pQ����������1��T0ya�{�k=������ ��3��G��C�Q�5#7�曞z�*�:-����+�`���0�2���RH^�0�>��Z2��,5��S(��Cۋ�P �ɡ���|�&�\�Ѳx[�fsb�N���r��i�1��d��v#�j�t"�X�;;��Ϥt���Ǭ�^w���W\`U�@l�]�Q;�^�\n�wd1��^[*�H�S���qR-�f���^yXc�b��|��$��(a<��>hi�c���o�	췴�'�]�����9�.��*��8�K� c��=�������x�'r�Һ��LvO&R^�T��_{����������G�U����vp����5Ń{������م��M�՞�۲�_�o����uT����.��BVm�<Gu�%����)�f��i�� ���3�7���>l������X}*�E�k���|��;��ݥx�8��Hz��<9�9���Q��\�ŞE�<2z_.���Q��;��r^��b�a�ֱ��E3�p�{V&�3Y��%���LڪfU􂸷'5�ACC��,ȸ5�g('�%i#A	�{:�}Xa��+��5:Y6 [��:��`��:X�5��/ҨNe�HW�5ȱ�9D�e_{�*��&�i�?��R�^�+�����K�C�:}��yK;��cP"v�>�d0 o8e�/ �%8��n��D$�pr�I����kf1�t�̿�H)+@���VZV�]>1]��h}�>~��ʉ���ԝ�JSb��68kC����XЊ|k��`D�F��Tvh�j"���#4�Y��>t)C)����8�k|�<��9/�!��:��T��y�g*A>���տ�B��N�"UQ:�+�\���6�h�)�NZ�Cq�j�V)�7=�ml�&����_��$yA+�g����nx��,)-�i���-�D���yDN1E�t��Mw�B�����q�����X���vB��a����
��J��s��L�g4�C�Oy�u#;`�9}�f@�`�a^:*	���6=���'�^4
t�,�u��`c���a��!N����{��ҹOe1d������Z����1	!� �J`�~�-���G���G�(�&6�:���!ʫ� �	XSb��T��tD��/��Y#��gexN��ٽ�]�
�B�j�!�*�0:�ӵ���6�����q��"�-���b�}�O&�o\�?��嗄č�n�ś�=�{���-�Vت7}zp�܀Ѝ�ȍ!���:�er��e[�9e�^��;�[�e�Q;J�Xp�ǳ��O�A��r.��$�s��Q`�uFs�o�H����Nd��5 �rK��^yn��#��'�w
�߻nC��.�ٰ���v�@K�H�o�Lo����
�,�%v2r�@~B��V�j��t��m�F�7���	)��e͸n�g9.J�w��0W����ts��2n���H?�Z�:F� �t�0�*��*�X�k��H@���x�a�i����&�Q`ey�&�����K��|�溝4��j�-	��(�*��5�\�g��[(���y���a���Z�تĝs�l*+�"�)´MPʄ,�vm_�.���e* �7��aUh�*��ź�AvYpd������q`��3떓����ES�m���R�f����R�s�sHa�)հ������9�R ���� 0�H4+5��6����׌���b<u[IԽ���e�94oyx	�S-�?��A�����;������m�(�[�S\lⓡ�׻���z�"���M��t�hT��B�ʰ��KiGX���o3��p�m$���9��8K_�p�cȤPC�a; y���eڨ\�QKE��-��q�(7T�ΤY�w���~�f�|�g� �?ARMPh��  6�:
�;�=^K�P]�V73i�
�X����������^���Q�馉�"V�����4A��;�n�s����WO�U��G3I	�I�I��g�� ʊn18�����h�b6��,�; X�R=���po�/o.��;��$��(��������3���ͿX�A�]ZF�Z��0\c2^@�S�	Շ���f0>}�F8�c�B��-'��fkL�ͯ��P��EK�F�Ǵ��!�Q�gR�+Q��uX/�%�:bQ�"B�VEou 
�2����Ӏ�O��?�$��0ub�4���#�?����F��}w�I�������(��Hi6H=�ic���Ϡ���)��<D8�wrJMє�0N ��2c�x�B\� y}�����<ԚtU�4&E�V�?�Od�k.�t9O�KՖ�X/M���`�̀lu����L~z��B����(��������Z��S\��;������PV5dc�^�,�Y���MuV�i��>�E�ubd��l�r}��f�4���c�h��I-�k(
�r�e�1|�,�Hq+�^@�։��O�@�M��g��f�Q�ZK+AP~xx+��9��L$x'��u�'g����W]�h�"w�h�'����N�(�è[��+	�nTTͿ����:�N�<�:9����E�r�9����Җ���.G�ݑ�,����2�_�nr�nG܏�
�DHj�]a+ή���}�>j��.�\h\�&6Ӕ,%���T�xݬ�U�W�.�������^Ǧ���Ʃ�"ٯ��)/W�u��������5/ijnϣ����o�ԕ���0
���wp%�����
\1ޕ�d�}� ��G{|VQ�%J�)_YeB�y ?�f�T�����%+��n��/<�z�J�ǖ$���?�\H�y�p�:����:D7�*8��1�}.o�3�3����
u��M&���UT�<�(=�G�����
Ե�c�w�K�-�{�;�������(��W';��Of���~�[�;��1�	�3��a�'vtJ�V�Va�>,`0�Y���)s|���@���<�s��[�}��"a݃B�O��o���:�yt���vr���2��/��[@�p�PU|�TJ��a|X��S���ތ�\�(���������b�*�(�z���6	MO'.i�b�#E�>���� ��E��ls�x(����D�z,��d��I�����,o����Z�U�9���@�AO3�O.
u�dmP8$f�b �`W��S�����ϻ����<�+��(I���(4�䕬�B['։7�	��;a�y���'�P����4���v>�WE�m�߷i;C���pR�&��)���I`K��
eJw�D�$E�.�"A����q�iA���6����е���٤���_��ы�`}�+��yo��J�� e��46�bR�=�c�b���}�'ʎ�Mܛ�i�+H�O{j�/S�3�Y��f�M6���(;��[���l�RL9�����+�~\�S�&a� �;�ۺ&����X�ӛȿ
N=��)��g�ew!Ԍ��ǹE�U)�]G�L'�	P#c��\���e��ntbxL7`F9L�+F�=�9�J�?%��N���'b�
���ۼ^����l�X$�k��e	�����\PɁ���i���b�)�9�C�uufW-0������<�EP+��c��hm��"U������� j�͆���j	,D�GM��܎+��B
��	f��X�{o�hv���ou�1����
���O[�<�M� �̕�"O��F*п�k�:_��P�:W�t��9,�a�TyU�l�W���=>�'o|�<0*,�NK4@?n����H_�hl���o-�m	?�n�<{t�-��H��8�9�U��m9载%jk��2���>��������?�H?�wK�)ڎ�\'�t�8�x4�Aُ}Ͷ��
�}�^SM�PrjaDϨ�X�8�Y+�y��(��-�2ф�S[J���b��������*�(��;[*��sb���Nศ�p��Т%jD[���;��!�/�dO�`S7~8�2�1��W���U��q�vÃ2�j��%�%w	��ה�R�����Zͪ>��\=RRr�C&7܂��(��Lm�&�듯F��Hf�
TZ�K"&�=L�����n[,��P?��c�g���(�a���=1����j���jq�}��-��6l��pa�ax���_�C覠:�R�����ܬ�G	�`;�e�@��>�����Ű�޵�r������Yˣ"�b�;��Y'���6��A�'uz�Y�l�fKp����.�}��/�jX5Cy�NQXE<sV�]�-��L@�-��-a %Rj=��e�e��W�@t]�T���d�\�Y�.=s7biN��ʤ�4Ê
{a��j�ؽ&	�.�M���3�g(��2�^������S��8��K�SDEH��W��#��Ŋ��*��K�4֝�����W�A) ��͢�v��U��ۯ��QO���18�vjZa<�6�(�����!�'�M�*�{�� U��riL˛^�Q���m���N:�J����: ��oR��C�>BY����e��[��i�P����,m/z(�?$��K�6�i4Z	۫�cv���)SW\5���<!esF���<�0LͤHjt�<�Q�w��;�"�Pi)����N�����6��}���X ���Җ�.!h�7��Κ����)  n怳/�b>�k�I�쳩�>9�PG���1* n�F����KC����3m-F���D���e�iɤ9���?~����V�|$��Jh[��P)�Ëw3{:��{��U_�>G�rĢ�#p�h�|���=|-�~������z:֯�����%u%�5k�lf�<AU+��4��~�a�f��%�}�oե��Ɲ#p�p�	�;%Ϳ~F��Ql9�=C]`�>/	��yC���lA�hl~l��wt��.������c\���Q���r�{1�^W�3=τ�E��a�_���2!Z�3�����8C�������s1R,
��F��ews�:5��p��L�rdt�?�0"D��x�=X��>�hlH����K��� � n�D��2�=7�|b���x�n�d �ּQR�f��@̾��Q6A4���Zh�*Q_��K�@q�q?г��M#\q��MY����ԟ�{���\{�2:(�j�H)���I��g�?k�8G&	�r]F�(��6�d�����YU��g����`����*h�C~yNKǗ]�A�zD����i���bF@$3|�xE��IO�x{���x��5e͈�y�+�#�v��8���e���r����V!�T��莓����MNbA
�����o
��tG@� ��	S�%�����f%˱Tk�N���&�k�:kO�j���`�յ�hd�M,*�%` &Si��H[�M�9��'7+�j�k��¼��ާ�jx�qJ�/&[�D=}�@a;Q0�5���	w��$ �3ߘ�׶lr'���MDP�`)�O�C�m3���$�Q˜ ��8�3��#�������4P�[M%��-�����P1s�my�G�����\��U��Q�eכ<��E�Nͦ�R-hb�*V����M	:!�rL{�FD)�m�ڔ[�ߍ�3��bIi��Pv����DË!�!@�ta�*�v����;�E�u8V���m�zK� ��
��F�M���2}Hs��bc���ұ�]/�ѫ���̚�5w��@)��e�Q䵾��!1���Ե���ln��f��<�vT��C�"R$�١�cZb�mU{��FMH��{"�ޑ��/\��b�����u=]/ˮ|h���di����$��f���uB������c]�{
YO<��(	"ET���k@��w��퍱h|���r⪌dlu�p1nE�2"�;�s����������&*h�_�IFc24#�Ԑ�V�jK#������'�<H;k�ۍ`�Y4�*�-t\���sd��'��ގ�q�B�H��.��p����үO�X��������1C�G+nC`� �\'�I!]�}���D��s�̅#�u �-%S���f����Zi-���L��A�j��F�['�{��Ԍ� �WS�GX#	w��s[��&�,ٽ�?w�r��~���bBʕN Z�B<��ʗ_��'���9V���V��h�.1aq��P1�g]��Dqg��P���L@i�eU�W	��"���ԇmg���?j��{%&�X+ʚZ�u��L矤�����������qw��mX/�X�+� �S �O�h�8���n΁K���䍆�K��u(Pz�Yxv�m�y��*�f�[�d#��믕� fn^3�RhB�'!�~z��� զ?�����10@Vx�$ѰIg�p���&uU��\EZ1�����n'�m|u(��˫Cx3g���bK+|/Ӄ ��y�ͩ3�4C�[Ȟ/Y-����&�Fwc��M�
Jb�H 4y��.�Zq%�t#��0T1���_D+�Zà�낅v����P5@ˈ�ᡫ�g���������_~��uE�d(�^I��{�����_�y �'j�RȒb;{�F��ՠb����!L�+��*��{}���\1�h6p�/�%"�Җ����L!n1�`�zS�����K�U�Un�o�?*��_f���K �l+E��b˜��XɌ:��H�V%4{p�VF	��s��Y���k��\�'����C6�Q#�|����Z��6��W��kt��Z���(�l��x,�o	�&kpQ���@�&��}N��/�c�!;��2�!Դ?����R��)�1.�&̅NN�S����z��Dc C#�H��0�5����Xe,����T

m�'O�	W�x�렆�#	3�]&4ARx�Cݍ�P��x����_L�s&y'��K~_��g��;�@W�Ҧ���x�E(���h�0Q�T٢���S�a �zK�!�~��/8�;Xޕ���|��R��U�F:�8�b/�t�G�r��9�Oƻ��������h`�%���V�6P�F�U_d�o�>}a!�3/���^	��
�]k-˖ �Ѷ~� ���,&��?���܆�۸Zu{<�5�=�OjU�؞!/���N��x�O喊>�/K��(1.C5�$�F�	��5��CT��/�/��͚i7K̓,IQ�G.\�:Xy(ʠ�u��T�	kB)&�ޢɬ�*�=�w�H��ˏ+Q�#AI3���h��f�������*5���x���1�u��dҫl=#u[<کH{F�w�r�ߝӸg�	#g`캴���Q�m��VapZU�z��"���j�qY�_�3���2�ӏYN:���i�+ϊ��Af�sС�����4��H�+���q��=���>$",��WV;�>͂Bg'�4��1�(�U�E�;��Z��" *
�Ԯ"/ O!B[�$Ŭ>�/m=�s0,�L�ɠ@�Îf�t�3���[�jI�g�]�$Cv<�/���׈��ݧ���&�gݗ��\ϐ�UMN��B}{��I�v�G"-_%�-���9����F�u,���鯶*iB����?��e��x��=�"�l��J��Da���5�E&"Ѝ���#<�B���Jz��]6�*q �(}3qI�勇�	I��Ok�(�j��k��0�y�0��n1�Y�&�'�:icc }uw�,`�z���;�BW
�W���E$-N���������?�/���Rn�F�-s��(@��l.��U�3����������4�ЄԨ�e]��\���6�w"5
@,��=�J%�n���t$Vכ	�o���$[ENrq[G�:\QÀ
����0yTK��i�;m$ZT�w���[�[����=x�M^#����4���"���2K�������K9�a'��[��_2|�l��(�e޺�r�B�h��j�:H��"`�b8 >�é������`�ºm-��m���y�z��x2m����<6,ȕ֌�O�m���_IM���@[R�-��Ip%`���WcȑK*�8���Ծ��$�G����Z�6����v�oS��s��-V+���
C_�:�i��N���o�@ZkP�q��IW�κ��P�E4N{)�p��^[��DH���ɘ���\��,3V_x���b����'i���.�׳r|7�W��<�����H>7.�.�N��N��o�8n�m��j�I����VX2j.	m�xauY}��
��8��?=�#F��^�RJʛp�X5/�|@[�mɱ�L�1�w�[�N�w����-�cÁj��`�<1�����������x`5ۍ^_|7��Y	�SV|'�|�^���1�Ӻv�T�Ô�S�( �)�|IH����w�U�T�<A<��5�,��X�0_M�
���x���zm��޳h��Z�3�&ܶ���*���]I�'���K잒�:�7���y���T7Ҵ������{��t;��1����&�ύ\��\|g�2��+��H��zj��a�w���Z��?�\�nU�c/r�z���.����,�~Ъ6�a��<�G��L�W\'*�+^�S��\���{����YC��1ʇm�����s=6L�H=�#�b�-�z&�篫j5�%�_,R�F���S�i� ��	�?z�1���O㠉�0Ô����`�J��X[���q'j;\4������F�d�{iwi��5-���l�/��
�Q4$��;;�̣F���WQ�o �r`LVoh7�%��<u�¹dט �ivZBLOqf�R4S�[.����z���3�L(ڎ�Q���dN��s!� W��Nڣ���þ7D��ƚS}����Ea��(�]燌��	I�<�u���ס��q�ʒZ�N�e���"����ΥV<Hj��?Y�YUa�v�[-���,��a�r4H�w�/�1p�T�i��"��gB[K��*�Hꭌಱx1���^������`z�%R˹	h㚋�G
G�7�|�A�e�?D�eV��b�������y�UJ%^T6��S�:;T�&W[9��{K�7�A��˵��Y��Kk�	�s��Ez�޼l����ϻOY��Z����z	YH_:��rw1{v��f�&���)|�{,;4�`{�(*%�1��7��Ώ�g񱎟e�pe#VV�zD���r�E'd��%��}��s� `/�"�de�[���d^���g�4be�D���萔�� �k>��@���qMm��ɯ �G4��Rs)?��-�,�@�y0P�#���Z��
X��r��_<Ͼ��yDTA���?�1ߋw��$�Ds/����]-�-�g?�Wv-'�*<*�ؖ
�;�y,Y��|[�������BT�[�U�H۸4�k%w���h���ȼ^��@��~WÞ�����vV �,ᑴDh\m�����_�����UQ�vne���,L5�6d�}$4�����s-sF�D��hL}���&^20҅na:�5�D��v�J����D��ȵ�9�ٻ�L4��Õ4��v�&��z��*-vPȝ<�Y1 agr�S��Q��5z���Y�Ը���doGN�2��ബ�u�y6 קO4v��:��/���6A�E$Z��� �*������Ǆ^rrj�}��[���k��EC_sd8֟� ��jȵ}߸u)�w����-V��vV�n| �%�B'�4�\#q�����?�.n����`fZ�1�'a�Ī���a���	3�
(z��KA:q~|c���Ef��W�`R��O�f��X������DIO�u7�}��о���&����Sٔ�|��c��\4u}�M��D�x	jn�܌V�I�s�u���E<;���4n l �R�d����f;2��D�+?O�ΰ�|ʁuɌ�]J�mT��v���0���vٸ�̀��?!r�j����qD�O��vk�	GU��K��w���J�:ҥݏ*J������帏|�Ym����z�G@�as��z�]kYL�G�������K,s���/��o�M�����M�2��gm��U��=�/l���Oa�|i�&�2���9!�$���}*�`2i{�X�6�b�7ip7	.Ef�(o�(���Yg�͇w��v^
�lg~��&C}E�W�g_A�q���b|h��s�#��\aNK\��|'l�r��yޕ��>����\�v_u��q�����q�66v�Ù{�>�Ѝo��_E��u'm����j(;�lǚn���z1���-L�@6�-��P��:_l�������*��Q��vu��h�a�v;Y�����!L������(��#�:S�"����W>��7��];�K�_��fRRA@��E��H�	ź��P�����e}Y?�qx� �l�2������/0�\0�������w��=�-���?�!n���D��Hk7��Le����sWs�(z&�λ�*% �d�*dNz&^�/h�q�m�����&z���G&�M�xN��rC	܎���R�m5����N�cT��P�`���<E��v%�.]���r��*���{�)t��X.O 1�����+�"J'�����v����h:%w:��>X@N?W �pb59a}}��{�e<ɗy�w�Q\��ʐBE�F����7�c��^~��~�$+���3b��}+ЙŊ񆱏ʞ�����OF��x#���R�p�V��j��k�7kX��[HA\<�\�iZ�]��?B���W����Z^D�=YH���v�|Z�	cڄ��γ�o���)SVٯe j*���3+������n�)�gP�DxH�%�7�k(t8b�=,�n,lh�%L�˅��X��kLʸۮ���3.DLNS߳M@O��3=��<�Q��ѯ33�X���Z�v�њw��`�x������܇�cu�
/o��G0��2�'hђ�r/4f���2��jS
����.|�W��7�J��]����W�4Y+;x��W�� �!��z��q�Iv&����ٟ$�6�W��NE7J�( �ְ@p���p�U�k�6�5�VYtOZF�;L�+�X��	��$$ 3�W�{�;v�?�fحҘ��v�EvS��4|�ɂ�oO������^�|�4�?܋��ӎ�%H�lT���$�6{�� �H�~����'|���/s� ��
J^h�d_z�2�1i��Nh��M]��;�����ڭJ�N��	Ɂc��Kv�RzJP2QbI�Z]×k��+�C�+EZ\_�vY����+���ǘw=�:�C}m�i7��ۮ���(���"�7�
ds���9$K�a�"-{&������i�ӪP�߅n�p���rI	�����n-,�7���DO�q�,�"�����p褝p���^w��P�,�\t���eq
��-B2�x���E����-N�Z���o�P�3$�i��Bc�H����=3���`�Q��&�
Pp�(��	8����|m��(��a+S��pIry$yI#<�����Gg����55����_ۄK��2=�$�S��V~��Ն�������OX�/���� vJ�BU�ʼk2a���5�b�ȶ]t.��f&���pj,S�=�Unz�f�/�P=���[���S�}ʏ��?fPRC	&��h�����Cx�rK!�)�5�j��ȝ������W6 ���$��3�Ŝ��#f���!D�~d7r�@]
tj �Vū"��滧Z��x�bLl��pvi��zU��NфJ���3H�J�E�h����՟a%~j�^�I���wEN	�������6Ǭ���;��#����m3v�$;��<v��<k�C~@��*YNLJ�xcd]*#QK]�jѴlޠ��"Wbl��he߰Y��T��Šp�2#�Ba���8�s�&��<J�����"��_H�$��F4/w��Z�G�&o%��fv��2��[p0�������ylp�R(�DZ�Z�^3���|�ןK�C+l`ɋ����LQJs=S5�����ʈ�9���J2�co@�܅n~�,�5���V��ޱ���Ho<�NYo98,�(�
�����?#xn��)=N���F�u�����vM��'{MK�F����9P���[�^��iy��u?�vd��q��1�3࣮�(��{���'y��-�"��?j��Ug��(tg�-��h��Cw��Qu�<����K�G�x~�D�N�)�{r<s]	�8.�Vz�?���ܯ!}+5��� +; �T��ʐ>�������A[��#;�8�i�r8ƨ�.�!�r�CIP�P�e|C 1�]R!�>��A]kj:J�Ή���ոVVE86t�,(LvM ����� �f��\�?�.d����X	~{�~���?u���'��2 �ďI�*]{�Gӵc����D��6�u*�vM�lz`�	��c� I^j����h��� �Ҥ����a"}ѩ���y��ߚ���\:<j�K����FF�~F�H)`��Wk	+|��S�;��|�A�r��!C�Ϩ��Vx��C�c.m���Sj7��I3��N�.M�6lB�t�/���"߇�`���!;�V��O�1/H�U�7�`�c:�2S%��C�5�Ś�$@��Ie��1���_t��p�;�0+	.�	�R;L���c��\p�U�AVs�Lni��Y�i�JQ�k�K�@*��vZ�Z1�r�ZkA�,P��KliF�V�Ql[�
�6煲�x�b�F��wbh;��|�����3oN�V���;5�~���\��?�!��]:�C{r�g]+�]�c
+00����qV}�6�ݏ�0y�6�4u���?�gUP���d㾤f�O}��� �X��'�E�v��S 2�6)��.���Y�whi\��wؐ�3)�YV&�.U�X'8a��Q�/���R�$�i���(�?�)8X;��:�����e~8j��^�}�
��^��	U��T�9ûzE���}=�ze!{��%\����+��*�����!N�9��T*���#>.��[t�rUK�/� �aֶ��/�]�X�~l�`w��U8��N%�-g���<�V�"7�·�����\�S9J+'3&���8 ���*v��+w�_�	nl|V�W�"(��H�W(��Q��z_H�gX�\�/��HƪV)?١i3��H�4���q�0;�5�J	����1�$l|)�	��v�n��riZ2��r���Fz򌋃�{W����8FN�j��(��X�Y��v�GՈ t���P��	ט.p�E�v}�}f(�T+I�>pL٫Ӹ�W��cb䴤Ys@���T;xդb� �����9�BZ�C�[��Ms�}
�;K�e��}5�gJh�]y'�J�o��q��/���?L��j���hc�ύ�4�o�|�u��Ed7W)G�"��A(���竌����P�-�"2����x�9	̗K��e�a�����|­��r�h�]��Qk�S�V�y��;�Ux�`���0Ŵ����#I�T�~��O�9��/QAUqlz9�T�|H�����Zz�B-�N�� _
.9B�j5p�&�W��}��QjU<�rٹO2����82����.�: ����m���7�A��YW8Bn�x%�G[����}�QE��N:�����`9��|����%�F�G��Z�y�cvd��Tg,Q;�S\��{�'7�P>K�5@j@� Q/������k>�<��w��ы�)�h��id9�C/7z+'�]�T���w��φ$��\f�2ٹK�e�L��)�%��z�6�ǶA*��LY�F�%W��6{$`;�	�5�̤������T�c�N�2k�]0�`�(�S#$���պ����8ZA�(�k�Hf �.A�eH��y���IY����ɢ -��\z�1X�MT\+P��]lH�SMF�.UB�3�����i��[���Wʭ���$$�&�.�C��N�t�$Iچ��?�HTZ0d�
NH��6-e>$���w5ih
��E���2�q���@��Mh�=��K�l�"�|VE-��5;��4=���?�6��W��Y� m�r��<�-cX��L�י�?�X ����i��u\�@NY���,L�9�z��2�8K�9/4�\�@��D13�*5�b�L���}wQ�r���BѢ�� P�6�LJՃ��1�cA�f}�B��"/0T�|8��t=�^K=�IV���?��"�6KX�Tr&�r�VҲ����'FI�Z��[*��}F꩝x�F�t�`��R��.Kw�ڜsZ�u� �4Z�j���RD6H�g6�]gX�Nj굋qLBV0�X����Տ{E���n���s�V!y;%�	���Qn��TA�wqɇd6#�p넲�\̓ )\	�9E�-�g��g�z����c�$SV`����#v+/��"o51��S��J��Oo�뛃Z�O�|�?� ď�if)�
Gx��]� �:��3Oe�� �/l�����*�@��]�0f�4O�e��ܹ�L��T�^(���H��@8[=ZRq�v?�6���K�z���.hirւ� ����ԕp߀�O3/l�������&H,�����.҈��V�qE	ѥ?�+ꡋ&�ܑw���:!-$��Yq�����&�]?ًD8�5+Dlfќ	���6����{���n'u1ӝ_��8�%em�Ҿ�y�J��._z�
�N�����d���Ι��r�݉��{Z����#������R�GR��,X,i��u 5+�%f�է�ǒ��w�FHp���4����f�5v����Z��yA��.���!��[���Βy=d0��RmFy���h���;fD2�g_���ox��D�B�L��X/[};�Oo�U�zO="�Z�D(.J��қ��e�Fg�b|�͈��+���V�s�k�3����TNLT�*�^Jx��y�XЭ���)Ԣ��f�lL�/�Labܾ���Z��-��~:FG��ά3<��נ�g6~��'G�{�L��x8x���"lT"g��}�ws�%��K`�2�x�e����>w}5J x�m�.��d���_g���d��B�ruxt����|m�Q0����q'-'�QG��������^���t�v�wB�,�i�~;
�S��C@������R��-�C�2���i@����p-�z���dj��֠m�ƭZG,�����n�V0O�r�Uʲ�$�÷��h���]�e��p�8�jI3��#�Cu��Tf7�;o\xp��0T����� �IԬ��K-�]�ܹ�!{;����#�/_��֟AiqT���\�x�0���rX-av� �_���	��I`)J�Z��?TP�f��/��/��Q�J��G��(w�?~U��#EZǨ���G�}q&[P�g���������Ї7I=�i����<�3[��6:��+�{2�?:�EC��Q�ZTLP���Zr�U����/W��}���EF}�]�DS�d�_U�I-`
 E�����"F���Wt�i�`��K���#����k��oo��l��<�2%*�|��������Ê���:�qq)���l\6� �;��3��{s(����g�D��P((�
��hm����9!�^o'��|RY�%`wוؓDr��@�5�4"ߖ��(�a�s�9B���!=�2(��ѿ���7cҖ�zǩS�|@]����ٺ	�wn�{���٫���!x�x�wl��YD3��Bm��~pe4��J�sU�_`���B�-�[e�u#q������U��<���ߘ���]T��7Ӊ�2.�&���0�h��{���E�z�]&��gWc��e5ʽ܈�N�+z�T�0�+�>κ8��\ߏ7�=�bs��kΉk�J���sd��Z�~�_�:�[du�F3ϞW��5\m�Υ>Ij�f��-���>��ab�"<��,7w���{�P
{8�#�c���0N"�%��|�6�+vj�b�2�i�.^�vXt���Y�4�l��=ǆ��h�GMK��B�.ҙ��t�ξI^2���b7��#YK���'(�c�W'䬀�&R�L�m H�B�)Gn��I����	o�$��6��تR�RpHF�s�i>F�<��s��A�@9x�Λf��aj���Q�s�T6��/�yo�s�;�~�X�ז���<�A*���z�HN�����ĺ"7��P1"|�>��Ӛ�|�t|#p�y0�V�7�ͮ���ڶy���X�#[�_�F��q'�
�3��X%5m�U����b7V�i<��eʿ������a�F9���G���k�F^hF*�%���vEA�۝�#�塧�U��}�R<���Y%�505�n�pX�z�g�$�v����4��ت�l�s"0��8��.�N�3 ��#���cc�(e#*I��NG�۱����!M���=w�Bf�D�}P��G���7�]V�4g�m:��}!�R@������^�n��^_�9 ��z�AE�R˦L�:ze�F6�Uĝl�*ĺz[a�[��ݘ`S'�4���� �k�0I���^�Op�<�lg0�%�߶��������S3�T�݄�%�D�Q���y����ן����)�A��Q6VU�x��z�cz�)�ܒ:�6g�饥��+��	�"p���c�Hڍ����`��-"w�ϓ�R�̮��u�c��ׂ���6?�F�#*!אVd�S�CE���n�r�lf-�]CY�Mt�:?:��d}�E�@S�!���1�-b�Y"��h*�=|1ʄ�V�ً�$�l�Ь�w�0�'ֆ���p;��m�خ쳗W��8��٘�4�i�U�2���3*���]]�9:ر�o �6p�k�6P^��k`�n��,L_E�,@��\���9kY�K5����a�����	��o��\��VW i��)��x'�P�e�� ��\�҄+���4Id��^Wq�(�B�~�+G�j13�v=!,T���}�##����jJ����O�+(��Xp���&�+�4m�^{g�PZ#8�E�C�����nm�ɗru�s�7��+�� m�3��u��C����^�w�7��:�o���yd{�*����k�|b}��+cv���`��v��X�08�4%S�U���ר,����U��j���Ȝ0(�H�=K�x4�M����~��k{٭39�zt�Q����H�Fxh,d�D�s�]�3q;����J��s鄪�; $���&�H�ӵڦ�~�01a��������Ho��da(����Py��py�����q�'f3��A0?�Q�
�"���.;n[��=\0�-��;5Z�Vh��&���!4|:^�A�����m��P*J��|���DgCF`� ���>c�;Ιo����p�R��u���Ð4���7W�	��7���������v� [��s�[e�V�}̶%$#XO�~�L��︋J�Gy�x��38�&�}�D�B�������Z���h�	δ �\}�V>�B����o�}�-���J��I/��+�DO�L��d�[�S��7��b��z��J��/_El^�!��(d�qT���Y��q۸�\'0?�G�Ϫ�9��C��+�#� tI�~�"���i��y?B|ґ3����-�4�� ,̂�����f�n~m��<F����������Y�H�2�ZCV/�7P���з'�k������Pm��������Ӗ�}���6M�`��tpv�q�	l�`\��gˉB�G�d4�2���ѷaC�,�O��_�\��������	����2��K1�X��SodH��u���-����D팃u�ٳM�|U�������D�,�i»~g����\�bk��}u� �ד�'�_I6��u�4]�Y#�z|V�@��lJ�Y4��*��G�9���'�g��^�Ʌ���8��:��Zv��nʾ���~',���=�!g�{�TCr�1ԑS@�m�A��	�������d+��@�����kt��8]X-�+�2}T�M����~!�{�#h�f���i�ჱ��A��r�z<{��l%�q	�C��8�A��І�3%�-���1��g�U�Շ�g�e�C`�E�f�(��i��$��9{Im����:��0����创�`0ع�&:x��<����f]C�"_	�������Ĭ����:�adTȘ���tj�Y+��M�9�2�.E�c�}�?�L�\ ��Ļ6��P�$�hݓ�oS�f�k�>�|8��`�N�ݽ��������2��ar�#�«���w|��V�+7�0jj��-�.N�b���%c�d��+�٦��^��٦i�Ct�UV�uC纤h��.��c�?�`P�K��TQ8��86�$�f����VIAr4 i����:���WT.�Г_ÒV�$�mުw���Q���##Hh=���z��I)��.*X��]�K,�b��Ǝ�yr
��2�YX>1�6k��c��������5��9df3����v����Q�RK���Mq"%/&��{��m�[x�LN�J]dL�J� ���1:\pz��<:��=��#xp ���V���>�
԰8���'�F;��'wz�Z�"��J�Q�"Q���FE����Z�e/���}���!�(�����K��";��"8�s	���u�y���Dt^����1k�y�/���1���zv��yY��NK�諩 5�(�(�iۅ�7��ʊ��V6�s�~L�S�Av�_�o���3""�"حw��浧��3��2ѡ�g�BUV���� ��I���u[x1dZ�� {��ɱ����)����
{4�7�SWd��=_�i>��*W�2����~zc�2���Wz�3��Ύm�!i������I���j�E�r���@���w��J�U����}h�����d�>��ɰ(H�h�}�����GAw+c�5��S)��UØO��i�o��[\<Uߦ�@"��xi1SH!4��Mz�4�j_���+a.aW��Bʁ��t���;�q��[iA��6P��``�X�G	z�4��w<�q�	s�K�ܨj�M�l���z��g��|0	�+�2�Z/
���/�<���&,«��3 ��W�ѽ��_�miFN%'
���	�u_�������9Խ:��!���b���FeP��@]Uz�8b/�}1f9�|ÑO�m:eg��G���%U XI�$U���lz�:aDY�������6&��ˁH���� P��)+/����gr���(�\�kO[���[�Z���
 ������׎\�@w�Ah��ꖋ�핧���5��!�oF�*D�����e!��#�~=#��^:ٍ�-�碦�o�{���Җ��-%:��@�`|!����7�7�
���&oSz� ����E*F��7]G��T��'�Ѝ9����!#�R��4��/�����wU"�Z�����TkE/�������<;�PԨ����H�w���jy���%�N~����^��/�ͱ�詌�k�ҐS	���)bu0	M�#*	A���������j���T_���k�k3��]v3_zr����+u G��U�ݹ��+#�D ߖ#Hg�;W3�s~ �K�6�Xh��<+]tfZ*(���F�]�,�|��9��(W�op���-5њ�����}Ĝ��"������J�V�Ur6���D��x�E\7�$F�-�|������@��%�.N!�2�A8�\�_<$��~����Ԭ��Q��*�>���ϟ�VN�h���V[,�B}ms�쪕Z�~C��VК}A�WAt[�3�^KW9��|�F|Z��)��4�t?��+�ij�Mb�z�!yw<�n����s�~�	��l�$��䛍Q�:��rx۵���(� -�*FmD�d`C��l�)*��hഩ��R	�E��u�Yxw��@�^FŚ��­YЋ�MY$$��_��=���!z@�b+V�N~���_�p����˕-?���B��\�%���^�oC�d��{eԤ\@FUw{�=N���qޭ{[h�	j�?�!Z����(R�������z7�룧�֏��?T %��OhiG��I"3�����Q��oi�0�S*Q�U?;����;ً,*���M��/�B�����̷q	J[�?2�Y�}!y`�|Un����k�#��G��nRF�"'h{��,N��A�i�._zZݣ<S��zgj�\`z��I疁�C��t䃚{��.�g���'Ϳ
9QP\�	 F��͹�b�}8�^�nR�&�4_Mx�p'~��,�A!n �Ǫ�h�d�N\95�d�\�@�"˗L�6�����yoh褙�ѿV�ҵq��XC荦B�F/��_T��]5�!�:��q4A�ƚf��M�FM�<=��S��eD��A�`9ng�ph�T���<OR}Cz�M����Lc=�Y%)$o��:�����ͅ�����)�&Us��l���jnt'b˹�\�E��و�ƘHMo.�z�h0^ ���#��M}L�-Ȥ�K-�rIZ��
�'���g�ے����������b:yw�=�� 79�\�����=1�'�ĘB]]��%���y�4r:Eġ����m5x�rh��OD��*���z`��ͽ?N�Ha0n���b�Ы�uy+�Vf�� ҏ�i� �)��s�2�dr�0���*��j:9JU����t��SL���vW�Б��%��Ѽ�R�\P�N�f�M�N����R���TPLp�Qh�e�g>�����s���6`(�q1��e��Ē��8 �Fi�;��������҅j��D s����u3�ֆn�slx��UӮ��|z�e�y�����$�Y��Z�Wy���fV6���&��zh�闼�˦�̬����PV,#
a�_�|)�e�ơ���/*��<�6˖�t%]!	DOT���t��m����I�ۆ���@@��8�O(�IO%�'��+[VsK6�"x���e�ũ{������6!N��WZm�J�M��V����ROS��<�Ss+ڎ�
�!���z�dY��8�p�b�"447%F���#�F�'o,Z������f$��g����9?� �Y�a.�l������΍����F�,24�����0=���4Y�:�0\?HGp5uN��_o�W�/7��F"�aUZhN����h����͇S�\m�ʗ���=\^�BC�P�g�(��U,`/m�W	��JҷX�zѦI�jQ���j���qzn�]�19S�Dv��G�GHP�))��!��:��P�'+ځ%�̎�R���%F�lq-�h��<n����p�i(��;���Z���ݚ}a(՜�u�j�R��{l�W��?�{�z�͸I��Ғ>�_���!f��ә��:�<�����3�gnB|��ټV�����#��[���U�����*��6S%{�ؾ܍�0Z��ݵ(Yf�O�^��i�z� �I�ݩl�e������f6�Ʌ�b�F�$�+>{�x��	ƍ<;c�a�c��C������F�#;Y(1��j�b�'|cee!"�B㮁P��Q�a�s������?���YR�[��{R��"gW�]���:N 0(K���S�e3]���s
i�'�A7�_d���D�Ԩ_���A�I�l�QH�gE��\�nH�VhK���č �����h~�H�iÐ �\����vW�_�d$?����va1��с������^k�> �͸	�͂�eϾ�ƈ�a��9�7��bn�N���WLD/��ui#ܝ��=�N�������(��eI�Hv6����c.����F��{�N�W��NeQ�a�z4�k]ޅnt��M��҉�.�����p��N&�<K�7��]ٯt�O6:�/l�˄#Mqo]E��^�g���%����}�oܬ� �&�;$-x�	�2�&����|�t4��އ�$�C��X�eF��/̥��ã������T\��lFI�c ˴�
YN�xh�c��"��s���ׅ3�*+X;�9�Ul�;-���CV_�ʈnN�cW6aS�0O�>K��I>��9rtꛡc��f(4���I���G����M�k�)ys��f��(qGV_ݫYAK8��T���W��0 }6?���m�[\���ŵ��Y�:���#Ե�FT۵?rv���yf«h��)�|�[BD1nݣev�b�[o��6�"q���#�ÅZ�J~���a}8�>����qJfH¡�zo�ءH��͗5��R;��Q�N��AB�He�d�О�s�+b$f��3Pe`QL��T���������
�F���C8I����-���B�G��كEi��o��%L���E��Q�	=^��Tl\ұ�q��fz���v�1�8h����b$f������ꜣBd�g&����*��ym�w�7)߿�5��A���a��ȩ�[���vC]����<��1�5��>�K�\ݲ�g������.��e��W�S#)1�p�e�? /�sq=�6
�vpnXP7y�GI�џ�QP����9 ���dC�.e ���p�������;�S9߼���c~Q�f9d����c������u�<���J(��~��\����M����������~7�Dݣ	~
��\cFhu$Nh4kΨ�	)��و�7�#0w-|DK�)���վ[�<�3�¢X���	�� O�-�W2G���3��oӧ��hA�^�k�=����`��y��gu�GyR9L M��\3{�?~E��O�srl���ދ��G��-�c5,��KUD0�T���#�\�<�ІB���|�=�5��!᩺=�����
,�>$��[;J��i�tH�9���b�3HkV::�ޠӧ�]gr���*�P��UN�_��E��EN��*4���Kv��Րġ����]��'/kg8��/Ӌi=��k,(���u��*y�) a�E�K����W�+d�e�V�����Dn���D��pbu�q�dI���Bm]���Xәy�c����w��+��"P7�R���[�|�Ǖ�9�@��hc޶f�!8��F� ����7�UtK/(��&1N��m���.4X��<܁i� eϫQ��y���L�4
�Ɵ��&�b�3T@J�Luz�p�#����0�t4�����o���6h� C��&FL�2ʋY�+�[g#�nh����7���</��9Iy��ßEw��V� ��6�$�i���M�bc�D8�ƭ��y���k<�ү��%k���pcl�ôAj��U���>��%���e���u2��k��(�Ѐ��4Q <"�A�)Wל%{ڨK^/W��x|��ҕw�� �,NK4��>�}%��q���-t��;�U*c걖_�=��6c���%?�{���j�����:�]9�}��cP��d�K(r��	�s��+I	�p@�#����L�Յ+ٻX�oϊ�a���+r�`J�
��Q�w��D[4��8����&Jl�c�jGO�si�dW�濉�x�7p���ztlx�g3yN�����!w�P���*��>�P�[Ku�hY�*-�6
nl�{�8���')31�2� F�&�t�¶����
�͔��&���k��@]��)�����Q�1�	�4R��������«+b=>�-�b-6!�G�Щ�Y����&��\���oۣA�C�e��r_
�;�O��2t^,�@�_���.w}�-}U<[��cȭNS`���|ݺ�/u|�t��X����v��itZ���y;p/��(N��z���\Y�':�O\3��w�zV�W��xQ/����9�ul?���|l������}g���UsN,2 )���qs�g����^@��@��'����sᩥ�h8M�埦㥓	e����5ِ]�p�6kɤ���Η�r��~t��.z�O����#�F�(������K�ZQW�|לC^�2��RA\��VK��aMl�V�
����1��ܬ9�E�*���C<ޣ\�Z,�hV@�	�B����!Q�n&��iG48I9���~BCY-P�}o��_
O�ǳtӇ�z�/��/����z�&��m����(�:b�I����5N}֨�3�1����,I�q��S��L�
:��['��ӿ���q+E��0��iS�Oxr��ߗ;DoU�=��Qg��h��	�xnN��r��l��{�ۺ��,>?��0q�.��L�Xu���供�U&�!L�ۼv�2K��F��5QP���!���/���=���/�7�CR��:c��?��e!��pw�h��s�d��%���k�
�H=kE]-4�]���6��������� [)��c@�(y�!BE�*hVl���Xp*��H�ο���Ȗ��������w��9=�)���PIAm��ݎ��_g�����)��XC�g�/_�"r���%� ���#�Z/����`�v�;�Nt��/D�l�u��N���T���-�C�f=nx���M�|�3�%{�J��Χ�|��.��#��kS��l�'1��vn%�t@,��>�+�[�{h�d8�_c��U0Y���n�7g1l%��}�C��s&�;D�R�	a�\T�(��ݍ���`�+~�X�Uev^#l�bx�qZW�����Zl�%�.\��|�iT�����,Y�z8�R�Z�\���a��=!��8%��*�|	4c����6����?-��&���Μ��KC��j�x%i�QoV���c�����r��-k��N�h��xК1<J�25\�B	r.���ޔ<ċ%.��T�/!IS�O˃K��a��&�c<1��k�Í��>I�	j3hF1��eۙO�	#{v�̨5���Z���@�p���;��i��,��4S���z�F��`��X�|��,���]�~�����W�=b�I��Q]s�������w)Al~�Ⱦ�W[ K�
��%7xWF>:�b˃ޒ2k�2�J'!�)�}��t��i���L�6{G����ɳt���y��mo6���w�'�sT*=Xn����~��yz ��kư��K6[~FL�$zE����ƵSHA3ldK�L��	��*H>�J��k�2��=��<#y�d�ӵ�3���!����*bUS_g!�lG�Gq�=��y���^�C�"��3�y�n��[�����SP�e�2 1ӛF�^ ���@��{��qrr6�2�5��uN�bV�M+�'�N�����j�	��N\�E�Nrn<Xq�IQ���*�n��'�5_"�?�G{^@(C���&K������#x�â�.��}p�r>N.;)|\�`�����_M���4x�T߂a���MP�<��l?g�Ǳf�M!�#�@������?{h}�.��%S/���E��ό�/���-���p���\���	B��: ��Db8�턃s+coH�W�N�d�܏��?�N����S�I)ȸ<�S��1���{P׆J���a(6�@�f��{x�{0n>��\,`���G�4�}"��Ǻh�f��'\'�Y�`�;��嶈8� 8�Y R�Y:J^��8;5���qH�I�n�(��#��:2R�{ԇ�ho(Ȓ�o��N��O�A���뀓�/ϐC��kS�-�����S�@3�oBQ�^($~�m>=M�l����چ(��+���0������b�'�NG�w�g�$���#�l���+��2�e������9ºՀ,�dx�t�5�Ԯ�2�Y0��Z��?"�pB�[�Թ[K�f��5΋�<8q-���r�f�q���ɜ��$|��#�\ї7����zO��&��5Pz�t
���TL�jԜu�,t��^���c�k����@Q�c<
��!���S	��1OV�Nz|G����L'o�S���	&(���ͅf�g���-�����^tFD�T}��b$�F-�x�?V�x�h�6���`;ĜfP�����Yr�;΂�]��t�N5��jm�ړ�A����=�Tk$l�_(��_�H�Tˑ}Y72���Z�
�oN��m�»�t��������ؾ`0�ď�����l����_ֶ�c��Eqx��&8�@��@N�	C�eؑ�ڍ����%�W�IqQ�F�|��_�ig3�Zy�o�̄$+R����͍�
�;))�/߇�HB�)�L�%.��TvY{��AU�F���M�������t����m�A�)��+���������t,m��S
3�Р�OL��M=6&�F�j8e$�uI�$
��'�5E�H�i��A'{�c�אsW^x�e9`{p{ byF�C�,�±���U��C�٦���>��QU�_.!f�G;��(���VA����;�{?�Yu��qN����z��3\@0��h��H����
o�-�>�JzNl/�I v(���F�w���7%�#0A����w�"W�5���Z3PY����5��(�}e0^��ڰ�!���c���"�f��&�x�v��@�u���'E�rGA��u- ]�
��S�c�r�0k@<B�+��sO>'�&�D�C4�P({t�����R�G��ᶽ��9��!/����y��Q� �>QWn:ޑ��!IJ�5ŀ03| ^{������Y6�;c��!�}�y�f��|ߖ	��^@����2�sr������nj�x�X[_�p��������5١l��Wo���#.��:�r���h�P�Y)���+����!ߒ�Uy�eyf�']B�a���ާ*�#m�p�6��Gh�Ӯ��0Ӓ���� ~!�'r9�!s�{=�-�UԪ�^�a���&H������G\�y���, ��Xl
���2���$U!y�+e�h�{�z��/sѮOIK�p��2F&,�P�Γ�Co���|�8���f��p��2+/���`ge�/4&�|�֊	v
���V��A.J��8+.eۣ��Ր�<kl|�z 1|HP&f2E�d��K�pO7n��Q�	�m2��W%�,�1Ⱦ7aj�Ƀh�Iط��� ���{��JĶEr�] +��pO�����z�tIƒʆ��*�`�k1�>A5R%�w9AF�������v
zG15ɤ�C��τ���q�����o�?�&.˓3;�?<�֨�8P��E^»>�!h`D#��Gx��g=[aQ�qu�d�VKY�k7��p(��w��D�"Y�WJ���W���*�k�榪�*����PCܰ����:u���,�'�3cE�Y���v����d�;`�0q6�N��>�e�� �h�^�t�,,�X�6�f�ApԾI�iǤ���h h�"�$)۟����! �Ƅ����Ի~�thf;�2�5�;)D�t짾�l�*�n-�t���̦��rD)|;(���o��;6�&p��� �>�@lM2g��G�4`�`��3�{�@Qv-�̽2���X&�+�7Z��(~K�^T���?���	��+ePj���x{ ?����l��:΂^�=ecc��_��ϔ��}<]���q�"]����-b�[@[9�4g-�4k׼����*~����\�*���ˉ5�U:-@������P��0�|/*B}�t����b�"N@�#���>;ΰ]��)���$w{|�@�������	��6M,�1I�C
��ϊ$�3����k��_�n�%O7�+�s�l�.����=��^�3�E����E'`i�t&|��\>�(���� �_u��G'_%� #�9���-������T��� ��`��2�uh5g�>} sg��+��TK�*S"�|��N��{$\�v	���Ҿ�k|/z����tc�Ga��+�F���I�z��n�L}�L�}�ӼZ��nT��v!���fm��8rr>�y�IE�����������>�5_�N��g�Qf�2�`�r��U�U�:~���D`
I�.N��F��[��}���JS�а��¬�8��b�fϼ䶧/�<�F{����np�p�/J�(���qלȹY-RI\����Br8����(˚/�'t��λ}o��]DĠ�L��R
xPQxJeQu�]�ِI��e �?�&�K�cj��;ج����<��)�7� u����v��:4������U,�<�����̎��
H;S��<�)bg_�'�8�2�
��\ó	i�Jw�gLE�Ӻ5e۫y��2�i^�E!`����z攫d�^H%��!s��������ɩ���H]F60��Y������y��E��V�4�eh��)��s4lh��K�w�;��f.⎦RKd�R�C�[�ƽ�GB&Q�@��dh0�@Z�~��G`F�*+���Xz�cd�����prY�`�.��E��`��nΞ'e�(�H�1��ը6T��}��� L@�T��Y.��F/��P�6*����­��o�)w~ �_��V��?x�؏�aM�O�͍��T�!y�D��q���0)oLp?~�)q�&�Dn�T�+����@�r���X��_�w�)��^�BD�oNM�!�r��&h�Z��h��ʏ
K[�Y,������9��~2��]�ñr�L�kդ"; �-�&�
�?�ϓ�4V���B����.k���*m��yLE-�uPp�T��;�]�iSz���2�KF���ʞ�o�x��CI��,������P���c��>/D��e'lwL�f"��=y���b���x�r���r\�_�r-�6���h�o�j	Q�O@ M�"�6���1p�����h:Ɨk(���1u��2��;[)�W ��������ɫHF�do.����o���C\"��D��O��	�%��d�|�R�;�d���cΓ�W�
@ӹ�&菀c�� �QqV�'���xL�!��V��řȧ�t����Sj�杣���"�R��j�������g>��y�S(��4TD���hf��Eoy��m+*��P���ּ�����~���G�������-�O����!߾�I��;��Gx 	���]������J���H�<a������_aS��͚��<z+|B�g��!u(����?G�Ê�[σL���bݤ�٥��_VD���)�:/�Vi�]+3��kӣBt��ϵ�D
�0�A�I¶:i��!�xt6�*���\*%4{�M�������1�4�Ƽ�o"�*��$GO)K3���D��������w�w�;љ�!~r���H�p���Zo$��3!)��H�OU;��&c�a�U���U!�P�ANh��L��ҿ�����-׶��h���d8�FS89�;VEt� Ws��0���X�Oj��Ќ3�Y���7]��2KF�?�=�
L-��Mo+J>w��'H-����rg˚t���u��^.|"�<A6���B�ky�ɲ����ւ+WI����!Јk��ӿ�D�Q҉���3�$�����p�z�_/Z|�T*XɈ]7|w�q�mW?���0�Ml��֗��<��O?y{�CJ)���pr�� ������NwD�v䪠�����+"t7D`I{d;�"f��T�R���=��x�&���ɮCa�Eq{��ܭ���]9e��&�����kI�4�n?؋�����Q~��&����M��w3���NV�+]�q/����O�����_{�����M�c����T�Һ����T0�4∮���;"�*V�Z���$�L>�͊,�=�{W�4���'7�5�*7
	�2�a����7���SjHM2�+���C|R����WK�l�Y�]��L�͝��M�d��!sr��Y+�
�9k���ϯ|:07%0�4&{��K�G�J�Kj��{���h[�U��`�.ұ8�����5ڐQk�0�d��4�M;-Մ����+ u�}����sβ!o^����O���dr�<Zi����Ʋ��^���qi�f'�ܐM���k�������,�m�p�d�o�<D���0��\������mcL)E����x=��`ֹ�	2�TF,#z�L���+�u�Q��у�x[���9�ʯWX93N���$3y��H�_1�ĵ��!��m��?�3�B�5��nu�jkC����-f5�m�$C0&<�v�̨��z^,AT�,���J�'�5�:X{uF���j���V�ۯ�H�"˷� ���⣇"po��������*"\y�c'J˶S[�[߮^����C`��UJXT��C����.��3jM�B7ts���o��7�����[3��L�Oֳ���]"��`on��;�Yp��e�u7�HX�P�`���NLZ�d��{�q��E�zIi]w�H���(�܀4Wri� -HƵ���g�,r(�H��l��R��C��I�}�W�c�� � ��Vʐ��>˞Tj9Ю,+9򠙘-�(�xF�� z�Гެ;C��"n�$v406���B�?2��b(`���6�`|;�#1�����bQ�U��΀����=��$�w��t�F7OM�e��
_��¢cX���8$P��es��j�<�ݣD�J��d\b!=P�&B�����^`2������1�g9�L&��'\���-f����1��r�R��,��Xmwjok'�ƛ�H@B���7��d|u��a���bV�\���TU���OH��y`�,"^�w,�wk�8�5��������͘�ܿ.-�dC�5f��YM�|�w���D�͉q-��s0��dFЉ;/b�&�'��x�������\��t�Q�o4��hw��c!� �F�r�z0�?h��轤aԣ2�;(��4:���SƜh$!0������JZܰD3Ss�P�Rw˴D���-�Stb�o1z�8��0=S�2!�[��X%l��=yA��L�}k�?0���{Ν	ޚ���pKd�酻W|~>��β�Ȃ=q;�_��ة��X)A�֐�!�x۫�`�k�U,��#z�e��k���g8���OK[>�����=3�&vz�&di�/0`�7%�ϫ�|~�Li��2�b�Ŷ+��A���.3��n~��-��w��@Z�N�e]'�Lc�;q��9�A5,	��"�VS���^t0���^����z"�yJ��7�tP�ZJ��m0�l:#��aY�ĐD�ʠ%���j�����h%J�2#�T(�Y!z�p��c���ݲ�J`7m(
SB�q#��i3�1��j�6��+.�R��8K�n�P{�C�Ӭ%Y�И*p�)�����6�:�gTB;�ݏ�e�2�!�*pf��Ɔ�Ɓu�W��2���<���[{����zۚ� �6?H��+)����VA/�'�`K�	���G�Цr�I�w���b2�]7�k%�[xI�^�� ��W%|M�<��`@�O�(��W��2E`��l{�Z�"��7��JZZ�'C������F�������=2�u�U���dW[��Hx��@l�K���O5�Y�#<=65M喴�8O�>rMcX���Fz�M�I�Y���{h�Jh����Jcd�����W��Nx@܅XK\�+m?���U��ІnM0j�` \����k���D>���D�~�xJ!��U���3��wb��^�K�zJ�m ]"������Z��#���OԮ���QO�8�k�rk3�:�� �X��2qp����˸���$W��"+Fuz��jb��= �883�n�w+���Kz� ��!��nhABƄ!(�Ψ�(�!鎖N�Va�D��M�t�c�5�.�Pn��,U��-�3/fo#��]}��	�S�X�5��8�-���p)�u�O�0Z��qݞ#��Z�=9� ZT��[%� ���ސU��.1����S�^#Ƒ�A��µ��}�ݱ4���l��u�*�I�x=ǌ��u6=t;
w":{f��2��|�8)g�$Ǌ^E�����v�]�*����ω:�/�p��k����졺*w�Ӻ*'��E��:�	�N6��8�v��:x`#2L���غ?^��i��B���XO�D��y8C}%���.�%����7�}!6�P	�h�)z	(�����Aύ4��@���~=�vRΟ*BS�s�l7q�A]t(���Fw�=��?���v�tF�U���i�)D	��������ٌP�-���iϖ`M
�����o�����v��Xz�!8�S���Y�6X�i�=S�T8Da�',���%��'��;
�:�>�EP��YY�c��E�C2�RD� ��}�b�8#��M������
����MbOϞ�U
ꀘ�;ReA���ް�h�����8m����
W����NO�h��;&�C���e]��p�To��Q�a�jx����՟�bp�S�Z�A2�� '��!�u$�p��~���a�c��(g����QnA��������9^�8Y>�1��`=�l�Qg���S�&�u�� �1}ͦW�ؤff�d��N���,��Z,JZf��C���]5��{�J����x%�*�g��ɬ$�<x������|YS�)̓*�];k�q�Z���c�y��So}��R�*�d���d�JͲ�.-b��̾j�����ݔ��E�ֳ!�X>������[^�Ţk�$/��h�������s���>R�
6f�Z�Vx��TOXc��&U�i�Qd�a�{8�� �[���ٟ�A�l]�ֳ�V�	9�9,g��/&���E�Ԓ��l��y�"�ȇ�/2
�8���^t�=����F@�6'���u�7�`0���5w�=%g���=H7�1;>b��]ـ �g�U��I����N64��L%*����M���Κ�К�;��'C ����=�����i���i#��U�I��fl���c��4_qh�]��O���fbU�h_)����"�P�����w�7�'�� >�pΘ��4�go��aoɴ�I�ۡ�JɎ�V�ą��NGt��K�t1�+�?xݸ4�.0��#��Ʉ��E��r��[�)��X�ֲd,���[ W�*��A�mou�0���S��'}AE��z����^h���3|�s����?
���3����R��"��l���� � t���~&�~�5px<�p�{1�(l=�yC���"�����[�\�7�u�{n��K�m
ã�Ք˪rʇ/�4��~�U�Z��5>���gL:�qI9b0�<fw�U˕Z��6��'V�[�����!5M�|�B��J�ٍa�7�;�����#n/E)�[��*á?�x2�m�KoV���Vu�؅{w��]�A-�[������;/Pp��H]O����mUD)�6�T������>�#��������tp��'�g�����ǝ�mփ��������{� J&q�z�wC[꨻q�|�MnΟ@�hdL��S��PAW�b`�)JG��hMB�N���gK�&R�ՀC|���yD�I�M7r�'���Z�J�c<9��)�Xا����`1y�Jg��妊�n1-�X�ri�к������x��߂V�Mܼ8$!��p��hkӪ+[S���`���Ά9�{��JCնx���c%�rO���U�5v�x��3�B?0We��ۉߎ�h����6�z�=�h��p]X�X3�E���[�;b�͌����p��#[�.Z(I���M���NJ���57	��'��-��[J"�3%�4��`��m�'_r��|no�A�aTR���wXR�l��+VSB�sQ�77=L���V��������󍚕%-*`���:I�V'��se%dDGC��T�l���b� ��y���~���&׏,�z�
fl�ĔpJW�������:¾M��:���� �G�u��8�q�7�`�I��8*B�0�]ٞZ��wm<�Pk�-
�U�L(	N��0�7`�I��$���&�0'`��ړ_�?�I��SAk���`���t����ͳL0)@ˠ�]�6mM�3��+H5ȶZMuc��?��?b%�j�r9�E`8�!x�s��Y��K��.&Y�Vp�l}�%B(���*<�J��#[� ���h��Yҿ��:)%��V�|3NҢ%�S�*&�a��RT���)���	�Wq�q$��>�T�(� 9d)$ջ3�����N����v���X`1P�sϦ�V��7�d ��;��9�	�Ի�z���W��-����;��OQ�ȋ���M���ٌ'�cW���=���8y�QP$��+=�wV�gk��+���ղ���}Q$��D��B���;�2i���D���-r����1Ù���Ԥ��.SX�n׽,��J�\�]�6��9M�v^
�=���p�K����)���=ѻ:<n���V�׿�$�Ye���'j��јl	���?�v�͚�"�Ck#���#�ʶ�~��Im�~���ظ�@��
��4�� �(��~�s��S�Ȝ��aȷ�nO���J6�E���� F-���#Ix���`�O�}\;I_1ܾ΢�<:��/�1�A�������M,T�^G�s-�pb��@ͨ"���J�/2p�q�9����,MbZ#c����Lz�-Z�U@���
��Z��|��4��UMV��L/`N�km]��&JזC�O�4��펭�e�3vs����&z!��t�v��~ BU�JP��]�3LWUǥ-�嗟|�/C!r�8`N�5���𚌣)3��L��^ma����p�?7l�e
���R�)��6#�X�T>�qи@�%�e��V����`Mxn1��T۝�nLا/�77C���$T
+ovG��XRv�w���#yf��{������� ����s���8-�{��f �F�H�~���
��;�r�߇}�|X��[>���OxaK�9
�?���g�sh	��~;򎻸E���)P�F1����-e���h��|�G/ɢƑ�QNҏ�s�(�N�a�7���f���E�ETV�0�y���;~}���9��Bw 2���������KMX� �|d����;q�����S�n��]���#"��@
���dQ�V,��#����:ܪ�����<\�:C;T-'B���H��z�+3��e$�P|�Z@&����Q�ͯ�w��w=N��?�B/�O� �Ƭ�Vj
>�����_�4����oz_����]��PM0��W-h߿�8�gk���B�|2_�]meK�����!
�� D�E�>]<����,��m,V�Fy#j��t%�=��cx٘�N&��-D�wQ�5]\�,�7��'4�����`�U�������ף��l	�ܰ��Ul&O�.F��r|uQ�Gt�S�f4�B�����;�O4���1/4b)�P�r����M	�N������M�]oZ�[o�(9�<�\�O�_�~��{�]�d$V��Yt��H�X�c�NhsY�q�&�E���+�%]���?0ڝ��j%�s�&���N���+�z�U�����Ծ�Fr5o�c6�-�#ԿPFu�AC����(%�����+�1��d���>4dh�	���o��]G9> � A�]$�9�ui%�.� ��L���U�`�{�!���<U6����o����0���/������9���U��+�1s&|y��U���P^9�Y�kZ�n��K��4�����
1�\i�֥y(��V)�T�,��@i�boteISz|TfY���G��#�;VDA�gC�b��ʓ���m(��,�F^��t`p�G���>ky�td[� �o��}#w���VMID��</����|L�rkV��b����ǉ��Zi�h���x(����a ����G`_9�8��x5�rAR>�%��F3�穬�$,"5�5F�(Ԋ�j�W�W���K��z�ģHF�3@��z���>�H���"�6�}���\Z����Σ��A�Ȱ�m��Rk	v�:1
p�#f����@~�q/�,�gb8�ץڈ3��ͤ����p�y�|:;9��ʅi��)�A���a�l	����g�5�����e"?�i���ΓZGz�����w� �T���45�z�����:��6�������J9r�W�2Sc� w����&T�G����ۄ���*ogb������	E���WYhp��[�	�=8)��s!.��.?�F�i�"�Ȁ��3v�d�m�	�������m��<��C�߱�r�z������N~n��J}���glFr��π�+r�=���񎼅Q�=��Ơ��9��8�?�x'�㟌߃�����p�9��OS������H �F��n�S2̔3�n��t�Q��Z�=&ݭeM��K��X����b=v��D�A
�@��Sb��lh?�/�Z���Isu�5_3I^�d$)W���c�xM�it�V�ϡ�=�/�.EϷ�(��
��l��i��EJ6'u�1ӷ��>��Fc��l��u��ϕx���S�(���]�*n�M��[�E�h~���
��:�·�t�䍅���K���;��T��}X�	�QfE��O�|���� �����,S#1�rێg�*����]�B?V/�$=�}����cٜ��m|�~i:������.� ^�k��О[q��D��6
�G(B�WW�W�*t�I��\����Ų�8��3%<���箹H�j_���*�� >gV'٩�n`|?+{��/�"=1��i��-J8�Ö�JSh#�3VƎn�� �'Ri����_&e��&,��thXKp!�P�
q�#��Q܊�-��S��:�Z��A;�w�̣+,:��2���.Y��Iƀ�$ೡ����n��{�k��7���H<�j̽XĦ�j����\�?#�����X��i�}���4̛�%�s����]�\�HK���M��ꌛ� m#9�r���J;M�gZ�(W�C �S.�H��Y������w�!� ��v�||3%�o?i�Y�p�r�����
{��̖i$`�<��9�$Q�6cD���	�k��x-r��Y�y�mv7���z���D�^1�%-LEI����I��X+�h�P��"7"�fx/�g��T��Z[+��w%@V�[ �.�:��B���,�rj	�2b�P6Ғ�����Ԃc!�#|ױ^ e������^���.�)4P8��v��z8���������� ��1Y@h.����:�'���50\�@�
d��c��2u����?�č��#q����K��Ui`��z~��BI���z+)4���Q�����!���_�*FSTh����U���tE�˥I��y�����"�P�B����_���^��G��@��'no��I�k}�W�,�!�
l�xp���z�M�m�6���҅9�y_,��+*�z�iʊ��Z�T��E��Bp�cG�2+݂`� �w�B�4�#U:-Y���?x����s-͙
�,��-��C޽F)��h/�,R���������M�=+�V#�Y�T�6�]��_ X�ɟĚ�S�3����8��;���Cxe�8���F�
�y�b�T��e��Ad�9�$��%EI�̧a���f9�D˅��dZ�`��tn"K�n�|�� +� �S3�����I,�{�h#�!,�6�g�)��_��V�=s�KayTa��b���)<;PP���9[d,����{�$|G�L��F8A=4
DI�r,F�\	b��H�V�2���{:�㓄� �Eu��{��)-e�)v�|�y0�E�U t�g���̷R*��+��O1�]x�w��]f�X���~CF� �t+�A@�H��U��9�"G������Lnz�n�aƛ�)�+�Qٯ����fڅ$���_�pz��"�*���N�r�T���2>�hf�J3��+	}�/[N(������- ����[��Z����׌Q�,��C�R�+�a{�U����oG����v�����{	������'u��nz;j�ő5KI��`&0��3k@���r�Oȴ���� �I��4(�L��Ua��Ej��T'�P�{��Gvt��Ԩ�gq��,U�[�����Ȳ��ً�$���]���YF��-ܶ�]Mɼ�4T������@I�	J�۫��t��P ��Ee9�G*�O�~�`��]w���K1��c�]�r6��v@W=Þ��`qEܒJҎ�+%Ϗ���i�o�	� �ntoO@�kߘ�9��QH�$�:�����7:�5�(��dt����1��d��W*m����AEr4:!���3�ǟ�U������:�J�����(���૸�`�y�9�tj��>e���M�Nf����pb�z%H� ad�iNڴcn[��T7�ĥ:��%��ux�N�jHL)�ѡ��htvI�z&�[�9:(j��#��JEmT��;�<�hl�ߥ!�ԷQ�a�Ζ�{�&���o����1��$��~.�K\��IFPRe�kz	Q$JSܸ����W:9�1k
�R�U4m58v�D>����am���p�2�'�_���oU�mn�N~�ʄ��5����,R9�`C�j9��)�\A*��P?�\fȅ����k���$�<:Q���2Zc+��ph�����i�>
0���$o��=w�jB���^v�#J��I�'�Ϙfy�̘d��f��Uj�����lƃ� 9gtT���qH �12Ce#�mӋ���&�4X�{���͔��� I�.�����c�3W;.�L���+b$�z����Ao9q1���[��קx;��0��Z"��_o��	����͍pw�������U,O篪4,�F�l��?�����PB�}��f�����%r��P���:ν�A(�pÞ�$��"ƟN�?���6�6�xm����ל�(OS6�a�?�䆈����3�,A��DD�A�6�0�ti#����k��K��� @��Q���~NZސشc�4d�/�~oI(�}�BXN�͗�(�;��Hk
�]\��ȨR�٭�����fD�W������b�S+��lH}�Q^�<)�)�$�#���?�ST���~�Ţ����
E�b�C��a�s���^I�}㚦-���O������E���Y��������G0�wS��㕖7�E�y��[���[V�@vk��1���o� {�T�ذ��r�����2�r����:k�J<@mW��a��!���6Z�RR(���,�a����r9a�|[�-���9u6�]6~�#}����ҟ��[ű�sW�jk7���S=��(&�p���Q���N&�6�$<~�)E�طGe3�ĕ�$T�5݋X;��Es�4���uA�o���K�XPO�<����Ӆq��B��y��~�2���襵}�c��X�pE>�X�:�1C�k�Lg��e�1�y(?��ҕ��G��{ަʃ��}ް�ZWvT�:�b�{����߷L��'��/]l%tB���Ja����)ľR ~t��m�QZ��6��0���g��/J�6�Q,���YjFBy�ᄳ��o����V)����()�����?�������X S��.ˤ�����#	l�ՌN�5�[�CGo]���|���h�6�\�ue���9M&���Q�[E��,�G�{A�qO)�����Ŝ�C̄v3�ʕN�G� @�%��� ؤf�rkuG^*"�N}��szA�z������M@��Y�4��Z��	�?;��+WY�I� c�Ͻ�G��"�wx|.N���f�y��1[,�`-E�m��Q�`fK����?�av��	�WN��Z��[|��A�1T���1���*u1����������O�ª_LR-��q��4��-�(9��FD� ��Dm���w��y�`eْ	�N�ɑ
���y����G_Z�'�("� wC:̌�}4�N#����{bh
Ӳm���刭ӳxW�^5O�d����D�B�����U�	�}��<C�^���Ci/�Z�'�H=˕�9[N��Nt���ԁ� �B�qn�/�?��}1�R"���3���X�_��G<��}ܚ���QjE����+�949�Gq���x���e�L��6��MU}l�;�M�4Y��'b"{?3���:w\e�N���H���p^��^z�VY�V�|<�-&��������x-���?��Y��G��o��[����޴�en�\��@h[ Ar�z�)��&��[X�QAlJC @'�=�=�'��>��g�!U�Y��:9 ���ns?v#�4~,���a�ζ�A1?		�5��O�+'+���Tn��)9PH�(��s���xS���f�vNc�F�i���%c./(�m�C�>�1�ɍ�x��B��M� �`��T�L&˜2%�32TI$�z�0�q�u�)m}a�����D\�ЄA�zf�1����~�)u�%�,�|u_�6���%T�z�];�s�]��~��*iFm�ԣ:�;�ru�g|��;���Mh2�IK
-$R47>�Q�9G�4K��Z�~�>=y����#��
�J�ɠF������p�?m���HlTjy( �)]k����9�B[�(z��җO)��wd��f�gX�j�|q)�����f�8�?A���F�w�8��	%G�	5گX��´�l��[�-��gJ�{�zueVR����|������'�Ec�8U&���]���Em�����i�B�Ip����*����b�z��W�o{�1X�v����p-�(�̣v�>�2H��N�o0��v咟1IX���t!F����S�Ûy%!�(�h��F���s�Y�+�,�w���C�
�d��g�p��߱`u�B;m����hT�����#8�����ȶqͰl��/�IX[-;�h]��>@�IN>ha�>J)4O���;���jc ��B7���*�y�p�N	Em�0z_��֪D?��{��uXo��յ�.����}��d
[���+��p�\hrB���*�>��*�yP�D�T�?)��w�瘎�S�`+A9	Z�� L���`[W�PF��7X|�������7�n��w�c�(쿵�����P����4���s�o*�FN��G�p���(�f'O$I��8J�0��9�&����q�l�À�+�*J���b�j<yn�2 �#�dDzNN�0�r�אk�v��u��HHsrT=p�a�
���e�FK�,,D��4!W�F͖�咙He4�D�4�s�Q=(ݎ���	]4Hdt.�r���Ȇ$5�~Qh{˹ �l�\��N�k{�Q�<`*PA5�/H��s(���*bP���4�Qǹ"�d_���I�͉�f2�pͪ��s�wDf��N��6�"�m���kt�z�\CӒ�����0?�:��V� л{�#t:_��t�`kH��A��Z��~��
jK$��5?Oq�QB�mR݇`��ka�GD께F���Aj�9��c����v�A��_�Vv�KCG�/G��,����P�OZ���l���0�}���S�4�#�"jK/~A�=��i(�r���tI��[u�-�r'���q8�CKC�*-�P~4�Ih3�,]R������Fd.E��8z\�Q�P!"�4]��m�#=	O�'y��^k&��� NOr�3�x��̜~�X|\������V?�f��P?��EZ6���A5y��Wg����ǀ�!fX'kG���Q�l�8��#V�#4�x�z�n�%[s���>�;3��\��{�����k^+�U����RY#��8ņj0>%�G`8�]w�?"��X�œ6�-�m�Q�Y���I�ǋ������Hc��i�U�Tݼ&E �.��@�L�T���;�����2"��(���C5�.�V�r����j��:��O$rJ8LK��(�-/C��bρW��,ܹ*�o�jQCC�=�1z�Yw��e<B�2���uO
}.��gA��@mF�i��Ѓ��(o���K���ݙ
4ޮl�l;1�%s|����J��Vp�v�36Se��-�@n|h|�����	n@͝G��T����e�g����<���od��\�*� g��˾}���@Ư��͑!�k�-t���HM7�l�
�T׍7�
����'y5�(�Hc�m���h��ӑr>�<K@ ��7�Y�b�K�9Xt�mF��V��W��ǩy��Cl��7O����?�K1�J��fo0D{��g�ڊ:��3��R؎f��w�w�_��h\�`���x�&a�0��$���l�#$0��\�§m�8|���3��� M����V{�nrt;���s�7G�Z�}W��i}�a������Y9�!����.?G7-5{�%p�M��ꯐ��|[1�y3�X�����ѧ _�Ȫ 2<aB�p�GV��Fnj늮�O�W3��_�d�.	�$6%����Z��0�LG����ǅ"m��J�2�~�Z���u^F�:�fE��hA��@�@��^Eer|�ٙ GzM�����jl��sT̰rY��O|!$7b»Hu]��	�b�-���]Rz��4M����?�+]��"C��CEZ?�=��o�&��Ve�!F�����A<���Cx���8Ey�ŉ��\~�z(x"j������ �lU�5�5�PL�Y��U�7�Q��Qn&,*c��랍�.W��+�+;����<�r̊��kab4,�{��/b-�]�°^~;ɱ>C\w�iK��HR7�TZ���^�5�0�}*�顗�>��Mi���h g�"lP��+6�|�X��G|���c��PI�1u���-z2������{���хxmp�Ϻ��ב����ut���*��٨�&�Y��3>D]��o��)w��@5����b�97�
�k~Wp��.��gH�nry��eי@�:�ت`z�jX=��8�f��7�T�!��u*�Q�K�Gr?p��at@�{�m�
P��MVkb՘YQZ^�e�7���d���������\�Z,�w��^\���K+aJw߁�3O�	�=	H�[�%_
^���=����k�mT�[r��Dh�DZ� |�U�1�O����t#QU�&+��E�\:V2�e;r�3`�����	̎�?�����f7�U�֫��ĭz�!.�N��D�0� ��e�|�͗�<��~2"Ȅa���
E8��燼Uƺh� P��}Hj�1�Lo���_ ,���+G����HJJcS�O5�~��)8zU �Y����ٲ'����tr��q*��Q�����Q��f�U<�<�\2�O#��I�\�|.S]JĴ��8�V)dmӂ�	�m_۷��y�z������/>��E~R���@ڽ�
�  �����)���R�����
	n�S�Kj?F+�X �9�hgQ��M`���l���ɍ���`�1ܕWTSOnZ�WC��E���q`,�J%'��q���o�?T����v�#��FJ���5�
� }�	?�C����9�VSʬ�6:�-��%�J0�	�6yӸ,��v^����x�V2�}<|t�=�*�x	�����>��혽8;��o����#Ҝ\���n㽩�W�'�U�o��f��N��	���r�p��^��v��*ӊ��A˭��S:����b�n״zB{�R�C��TF���=��_ik����	�a�>�w�H|���(��T��5�Im���+��q�	���=���Ꜹ���e���g�Q� q��c�41�4+v�����;X6�� U12�UuJn���6Ay"�o�0����Cu?�L��@������T�L5�?&��T!/=�@��!.��M���t|��0��S���F���J�4BR����R�EX�S��&V��r�F�|¦=n<p5�1��^JU{�S-©��{���zC16�ȡ������c�)S�Z�N����'^���pL�$���ؼ��6hI=�)��vl�1�ɵ����n�b�Д�y����04C�|Eb��5�q�;ZJ�^��L�o�3U�\�"c���[�����\�	%Ҧ�����%�F�E/��P���Mj^�Fu�S	������`˭r�����+���l��>e%�س *<a��#ZݧU��E�%/�'��W��O��I;o���\���L8���Y){KuFO�+������<>
S�Ú�)��N�\&��+\�*.�?]	\t/f�� >�F���̈́�/ �^C?K	�=?�t��?�K�l��,m88�C��6�aiy�]�A��pi�y�dB�ī+�&�b����vX����d��E��.7��s�E�%�^E!�G1ɍ�`��d-7��h��]TJg��r@bMGiT�>K9%-��1�&�@�.���U�;���a��`�d�Mځ$5 {������n��6��?�`_�N�;��PU��%�őb�9Wf�s��(k�6���7l�!���@A�<[���D;��) J<�2
�Z�T��6q�q�q�8[ ��]H��^zǄ?����#}�;"�@�V5�Cπl�~,�?����j5�k�pY��C?̈��|�ȡBiv��o�B)�r��'"k��ȗ{+��z�S�����U�j4����yQ�~�B�D�!������^�z{|�`�v� ��1�4`�PC��n�PF���$T��k�z#�R4�K*>�Pqe��5U+�����K�j�n��[���5ʞ@��S0X�-�9�u�V��O�D�77�E�r�:��.�Hd�ġ�l���aF�6���M�cmgЊ���!q�����J�;?Y��:�$��w��Cl
�r�4P�[��ʱY<����v�ˉ�>7����0���A���ܝ��[ԙ_/,����۳Kfj$s��\����g�9��M),���3x���%,]~�y��|��j�D�4)ΔP��J�湕�}��q..�vh�0�d;i̓�>�u���1�{�M����FL�u����a���Ͱ������n���f�|+ٓ����A�J��yv�
��W'N�b�9¼�S��� ������R�=o����ӎl1o~gt���\o��]�X��f>�nk��b���^&�ז�@�'�͆��|�e�S�h�	�����u^���La^��o��ӂ|���I`8��{T4IT��
�w������r>�M��(���!�dK�?�@�E��2͎�\�7�T។4bs�a��6�O 
�~G_����C/�b�5ϩ8w�E�7E�����p�#���էo��\����Ɣ���D9��yU������ۛ�G1�:�B�m=�M�Á�����U�����<ɮ����A|��ލ������^���U�`�c!~�7��Ғ\<;��1��t���lʓb.k�G�� ����z; �h
{�~��n���3b@�4)�hǁ�!I����V��X"QlM��{�kH� ��|����0���R��b��9���HR� ���|���n{����C�������-������0yʖd������ce�uP(���sŮ&��7�\��Vm���`�K5�.I�D@���q�N����9�� Uu���:3�범[~� �T�C���D7$B�ԉ-�E�é��/[Bf�����v�?�R��V𝚖>%䔚�i	��,��NV<=�?Sh%����R���qq��ܮ��֓��Z��ĈlHo��,��A^55%�[7�{$��*WGџ'���M1"�2G�wn��Go������L�o7�'@j�$ѻ�w�~P�]�)^����'��J�mz������e�o�/�T��0!���g����.	T��ٷ��;$���H?���p����D6���i�����7`plzcS_I����/�BGs���ұ֧�^��2s��m�5Iפ�Q<��-	�h�
�b%T���H�T��w��> �9��7���g�����uv�4E�2�6�����6
�[�\X�;�'��S-x�Y�5Y�Tvn<(q�$+�$�fR�`:Y�ǝ_0(
m'�E0���I�>Fk���xs�X�zT~)���9��f�"YZx�b*���zQjW��)*�Eh
W����h��h0��<��c!X?؀
XkX8�b�2
����Ŷ�v�Qܽ R�'�����^>q�T��.���N-�@忄�(J+m6�'5���/�'e	?{oo�F��`��H�W��8RQyQ�|2�dU]T�^߯=y�Q�����	���	n�c����8�r��8���6��\MC�k ��O'w)'�
=����f��[#չU|�̩����}�	c��2��՘Ӄ �m���:B$Oߛ`p���d"��([�$�,pl�*!+� �U��%O�N5�b����͠���Ӿ�fX{ŪC2��� ��z,)޻��9}��	g+��}5䖴I���ާM�/d�;�>��]Z�a�&�q2�v�\���\>�3ٴ��
t%F�����7�1�����e��!��<�po$()�+n�)�#,�ڑӘR�g��W�4a������jӳ`��}���lE7	s����K���;����<�܂X��$�E�{�����Le?�\8u*�b	�e���P��e�L�(��{,�'��8?����o�_6(\?�pH<��!��B&F[����a��N9�o[�wB1��F�ˋ]��%����h���#�t��w�y�e���������5$�r��D���-z�E+����<���y�}�[��sA�ݯO����;xs�DKпJ��:�$ l�M8�^J �,����ʖ���9?<"��i�pN��L�KR�*\�QR\]���d���wO[a������=sd/��k�,tL�r�vS�O�������{L@z��"����%��X�u��M�7B�BYN(d�O���\�&']�ⴴ�b���p��{��_p��.]�č�Z���`e�`��j���N1���dx'�T6w���>�]z���[������ƛ,���v�Yv�T�Ÿ���z�9�2�}���uf���f"�z	#�����%<>�4��iA�NI���#���?��-h��j@�D��ݭ����ݎ�(gH��3x�����E����Y��HM�[����Um�`���	0Q�nH����\���A9p�DR ?{��N�c�a7��[��PP	��Pb�3�>��_F��j}S� �g���n'<�E��$�)�G`\*-؏fH0����ԉ�*��|���a�-j^YZ֛���[��?��t?��x8:�-�'E*
�v�����r�X���CL�ZZ�Þ$DD��j��YyP����� r�u���PӺj����bI{�'��H)�0d�(5~�'����,4LGR�������AI�r���'�x���j8
�Y@=7���j�e�'q����j��/\�L��Oq������X[���Bۘ ��H&ӹa�ނ�
����'R"ϘUO�$��n ��25�}����!�ԛvAC��*Z�Y���g(�i{,쐋�u������3���fӻ�l&O���v56i�,��v����vR��gg��$�F�z�©9Z"SmK���nAH=zX��D��I�he�7�8`v�f/�$	�hn���n��X���c���Yr4@?���~�q����Gt���f{3��x�r�v#e�I�y/�]!m���1u���3��o�Rdjr����7{6�W���[���h���Z\�YS�ؙS��Ȃ}!�6�0#�^�b��2~��p/�(H��~&oj�ʌ�n�րj~O[����B��/�gԂo'�)��3�Aw޻@8@��ER�k�Ԙ?P�1�8Rՙ��&`!�@��:��'��;-��秼Nҿ����Ξ�Q��)�y�����h	.��¦�.���!�;4���tH�$<�[�����J�5e��&S<N���aa~%j6�E7��2/���,�Y�C1���2�4��tU��ًmb�������_�P~����
��%EY!�`)�
@��#�'�h�EzV��`���v<�9�$J�L}&(z�cw�z�:��C6e��)u/qy�d�-�T�-�F�E�y�:�����>דڵ�;5�?R�?K �`Dl�nq���-?ƛ�_�e�$���&�B�%�k߽�Nr�*8���:���|��ðx�T7�ֲ�%��b�����鮐:���������c#����(��N[%��7����D[m�4�JA�Fk,R�W����[��6��ZX�x����o2lǒ͟�������0@�]%@���l�׬_����ߵ�[<,G"�Kʷ}��h 4R�S�y�w�����D��F5�8����5�P,Ei���i-e��Q!{�Ր2���=��o�.8��
��ovIi���!��m�ھ}�m��Â�ٵ�;#=?�@ ��E��L+�"��(�s��1D&<�A�
�]�,:�޸ �XO�S�y��\�� �xC��H������h��}�C�G;bJ8޹'��!��	1�rA�m_x��4�|��x�T��:�#oW�u6�L�5�T2��O��+�1���Sc|�Ί�s��h�J�3��*�fd��-|A�gv	��3�%;� ��s�B�)���\\��ho$�V��mF(\�0�g�x@a����6�g��*��~a�E���������Z��%�W�N������� �ށ��p{�8�hP]�
o�|B�1n�xf`��!v'��{К��1�K�W}uRF�c��H�!� ��n�{sa$i��@�c�|��dD�@K�bI'o(}�'ڼ��Hj6��.�
=8����7kMi�$�ʃ�<�x���ș�yˏ+������$���C���5@��P�%p�-�<�G����fٝ޷�g����k��}��C���=�������OŶ��� �a����Q��i\]X���l2�H�@.�jz��	e�����yCtǩ.\pY�2=�7Ԧ��[��mh�����u��1�"=-��T��g���l56>�f��L�7�G$yຌ������|�n�@V#�Ʀ,hI`�����Uʢ`_���4���>��JӉb�9��o����cF'?��el�n�X�<P(D������,�}���c6�r%��nm������K��o��d0�/��1.#2��+L9�s�I>�}��>����#6���gUB9�F��%U�kT@�w���%{��&e�p�h��\D���n�<�_�p<����}�>��|m��P.�B���hn�_�CNł�g�&$�E
KІ���r�o�Z�����Y`>��GX	+��;o��fc����w���%\f]�N��1�������5��\]��h�_����G�pҞ�ne|m�D +!�GAZ��]�h�yܛ�t��t�÷(�U�c�lN�	�C�D���f�(ѴG�����������̑S����<v�q?ձ��差�r/eM���Ԕ�ֆШ�J�﵏��wԫ��rܵ-)�\G���E��ku*yW'Gn"�)�Ք��)j�<	����K�b湺����hby�J|(���wf��h�\D4G|t[�Y7���KMˈ������T���xޙ	��6�2p�g��
��]v��$�\�^��!��62�47����+�EhC�@�?-0ՠ8KQ��^.��vX+N��k&�p���u��D�om��Q��_��K?��/��8��A�t��(�w��+���x6�6��b�<����o�|rg������y�Q/�'g�.�E}��6k��cf�Q�R���mhÖ�N�
	Az�����J)�ֿs���
������U�;�h�0�Hc����Ը��`�]0Tu��7�P��܍�[�M��&�Y�R�Ɖ�_I�+Ï �ox�����<R F�:+HCCg4�.�v���`�j�Ͽ<c�%�bdj|��gv���[jJ�9U�7�H�s~�+���TL]���0I��E1��X�WjTW?�E�fwoP�*��+Ë��7�&�1�I^ �a�~;�șƊ�ǫc
�2���?�P�������+_ex.][�\�R[�-�ް�J�+�e}��w
ҩ�1�f��I�u�������fc�M�^����-&��b��>�s�:J�m�jon��SM����}|��e������h5d�%�����f>Q+]�e�
�� V�ȳ+Kb�&�b��F��>żu^vE|��5��� ��uZ�Տ`r$R>��!����	�F��VI��������0Du
s�m���Wȃ{�����7��̘�Բ� |V� �>W��jA� �q�yΰh\��Y�<n�9���S±i�GK�E=����g����b�GlO"�x���*ᒣ�Gn.���R����1ViYt�s�P\.̿n ���7�_W��
�A'L�"F��m��������V0���mB�6f��G9���N��e��e�S�%cT�A���Tm��v�Ξ���)�p!��x�i��0�ƿ�͗�;V���>Խ^���r���[�<����E���ɪ����u��X2������K0���6G�Є�4fX3��6�w�X�х���xP��,�p�k�P�XMS�_���������)��ms��l6s�du�+�8oIQ,aG�Y��Jm)xZN��D�1J�YY���kcsU2S�{~�e���ۣ��:
՗��U� ����~d"g�>���|�1��C�0d�)L�o�K�3�\$f��q�m���G9��6�KET91.�yD�l�{���f�<� �ǯU^�b����޼38a���<,'u�� a��k"B��$��?d���s#ኾ"E2���0�nO�a�t��jv���&��!a���>WVƍ�a܋�#����O��v ����ID)֗�L�A���Q�钠�ߛ�U&u6�Д�k�����]�>y����&�y��G+}hG����=?���@w-RB:[u�t�-�2-�V�A��R��|0�q!:R��A���2�ϘK�(�]T�r"�*o鄣�L6[A'�(-�1��^d��z��s�u�4G]jOT�����!=�?H6�e����t���;pFTN�d��>�jtզ⅂U�jB��|� �h��1�|6�n�fAc̒D��]�=k�	���C*<�l�4�}i%~7 ��ˎ2�p2��&3�RI5�~���#p�(?T0����S���"������#5�_{B��*�����o&�)�X}5	V�"TS0@�%J��� ~�n�B�3s�!8��/0�Hn��j�<�������`\��Q�	v��'��x�=g�W��=��v8nIpl����D|�͆3�4t/kW3�l��$&��q ܩہ^k���w,�w�:��n��O�E�����o5|�bw*����C}�����t�ہ)��y���\��n3�>=�
�\xS���Ą�l�yeLDh�5܎�q�Ze��b��S�H\(#��"�zK#���R����<��}LJM����Иm��N�](�s�v�3C����^�0.�]̖��;l/O��Q��g�M��_�����j���rmZ)��CΎ������$p�Hzd���f��֣q���%�4���opo�W+S�Fi������ٔ�:��H{:%��,�'��'B%�u�����JA�WT����"Cӧ��=�P��3�	[%U�?{��i�qJF�MHŐg��f��CP�>.�a,�Ň�U��ܛ_22�tvRp b.���Jȭ;�sT_�uӍ��,$sYl ��nc�3U�c_J�Q���/�h�>ͩ8S@n'1�Z��͉>x	�]m�Z9	#��/��F�K����#��g��\H�Y��'}����ƶ��6��4����%Ak��i;$���Ef�H�o%;]�$w���@�����O�A����zl������uK�f��	�P�r5�A��$�[$�ؠ�b�|�.rX�SF��un�T^��Cf;�X�o�3X؇��w�`zUgc���G:���T�m�^+��.J�)�ZڐQi���K���/�\�L�]F�FB]w�x$�����Ow����I�aĀ�P���֟�=���f7��lRyb�W��y�������W��Px��Xum{@y\;u@�����E�'!E0`L~NasN����7��nK���?p"�h�o�{xE%f�5ѓ�8F�9������A-�i�÷I��85�ڡ)?�A���(��2�;�]��u�~r���CasH���t�9E�)T�/��O���M��R~���ф�K��Z�)$��M����L1Sv��� ;�����Z��U9��W!�6��dRқ��v@�zV�s��9����:�������=�kß~���0�?ֿ����[UQ��|O�"��j�GhL���'���{)7���^�4�o��sL�|w��a����c�3w;����:>�$�i��
�@�p٠ؐ��!�p��:t�Ҁ�Ŷ���~H���A�-Rvͭ{>7~B#�쑜�ӂ�'�]I���|��8�~�S��y"=$Ȧ��RJ���rO�F�5���߱�nG/����o���,���O�-D\�p�t�7[g��C�۞WT�⾜��y�Y����X��k	|Cm���Z*D�����2l�����=�t2h�Jp��`l��(V.�u��4ŧ-�\ϸ���H�2&v��߻Z�!FΙsF(�Vk˽������c���Di��g�j�N�x´
��/[�@Y�Ζ0{����U�����0��!�P�>j�����Z��t�UK��pO��CphJ؛�'�$}�[��Qi �z�i��a?�](u[N����Ũ���)�20(��=[@Z�;�'���C���BB�o�I{"��ai��N(�E�6��[��ƓQ�
��W�xi9Z�:�������,I���¿��O������3� wt�$ٸ���QP��(6�w�9<US��J�)��o�2d��EH���8 KT���t}�#n�'�o��*����i���H�J/��[���m�3�丿��{#��	��M<�6W�N0�B>İ�����(U�e����K
M��B�T3䜳?���Ӝ՞MX��HΗ˔�-n��p�$�[�N�A������W�/�=9x��-�ES��m=C��Ό��]�}�C'ۿ_��&$�]c��9v������l�v��n*�����03-����)����;��BnF��6>�]��i�9%k������6$q�>zJ�G�4���X�Ft�/;�P��WP�O{��E\2�Xx`�%ߌI_�G�|��ܘvdT��5���Ӭ{լ ��I���UꙚ��[P�ҮhJ�8D�v~n�TP!�s��V��j�\n�������b=���9��cs�'BO�(�b=�!���8�\��1�%�R��TXR1��X���nY.X���f2�%���-�9���,���i� ���e����w�2�'���Y���n~�]w
��}�;����hr�x�V�Y���d�(�"ue�.�>�u?���m�td���C�mZ��f���t��(�*�Ƴ2"�YD��I=5f1�YfYR'(A�Y�I�}�YF)�IGr��i�s���H������i@x��F3����|߷E�i�+�.jL�}�Sb��z]���G��PY��c������:1IC���B����T�9(�"|�0AIw�ߤ�	]�� �vSSn��(!ke6\��[�����44�VJ�>c�����Z�WĐ_U
�`�����c���#fi�����t��N���ơ2댮�W��W�k	_ߖ���>�{�~Y����b��xI�+^J�	�+��KjO/���eGDǌ����QZ��kz�I��H����g�ݯ-��H�����;�����(㟃<4"�,\��xNat��\Q��Հ��c+�J0�{�����b+$�=�HTV�n^Vt˖�	���Oq��2��.s�Õ��+��?T7*�y�%tVɏm�0&����R9'C�J��[/��=d��Ћv�o����koen�Tȳ�����AC�7djY��������dfj&��OОŷ��FVht��72[
<|"�V���H��!��,3{wi{��]�-ciKSԞ�ᛎjb�Wͪ�	PzH�Ծ��N|�3�>c��&x)xZF�@8&)zɱ��*+@�>I$nh0�O2��#[��50_�����yG�7R|Iॐ�36H$�Pcf�d�����i`q��2�jw�mk� �Kġ.�8T����ף��Ƀ���գ����7��<ԩ�X���'��4݃�]�����>D￩�ǌ�a�X���@��&�'��j���a��|f�чZ�{�<�A���\\��u���@�A�E��tLE@g2�G���dvEsޙ���߯ҽ��@��#NȼK*(�F�؇��d������9���S,@塛�YaZ|Q ���?��m���r\�k�AC4�FQ��D_�M��TM�2o��@������J�)�i�S+Mdy-o��F��ݨ��N(��(|��'=j+��|9�.�X�2�,K�PU��%����wlv�i"��H�k��~i�?�Ϯ������V�ʮ�E�!+��W����P:HSW��8�Lk�ہ�Ѥ�];Ro]�s[�Cζ䳪u�9����=�TH	�F�P�"�!��1Y�(B�4�bަ=!n+S�{�o�J�(lk�*$�K�x<w]}��;F�L�g�K#�� ��sz�kg��&6tT�jmw�c��[����E��6$.j����}�©�ݐ�gy�$Xy�3����N�9�����U����t;�y�_]b7Z���:�|=�\�|
\T<��/���ޞD(�Ts�6��B�� ����S���0!wL�>Q�ҽ�(0Z[���#MN	�t;�ܙ�0a�@��|��w����)̖��)1U�
��_@ag�QY�������&Pd�֏i�0��-j@�
�j�x��O��
�9�5�E�|����F���>qiI� ~R~��iW��\�̍S�g�2�L'�񴶲(�@e�,Q�٣���>���i�s��j2���o���0f����5�h��#�p�U�_�[������?�@N�vZ�����Na�w��j�)Dl�g�u
��O�6�cҸ�O2�ӡ~4��/����_	��gt�^t������J�f���UH�V]��[|���Ǭ+�^��GO�����BV�����t�㵢�/��K%ְ�x��*yD3����#���gk��xDb!��AS� jG8�';̝d&Qy���ߤN�oK�bӭ5ԗb5;4�Ϋ-��I�&��Mܜ��8Y���~k������OD���&�B�z��J�c�P {0W��Li�(��Fz>7��-��=��=�6;XF����[1� ƨ��-'����m�:\����R��5	ɷ؀S�����@[�S������p~��#p+�����d�^'E�-��iT�%�n��j�_�o�5i����fE���Ú�G�՟kELnl�[�}_���X+ˍ�u����������#���G�q՞�9H*�r$�W�<T��h��#�'��s�ÊN�5����v#�Q���V����%�y�����D
 ��ZDj���{�\�K� �F�\�$���C��B*4�����0�ٶ�,�T�I8$ۂx(,��۵�JIq(4#RKHc�����5�0+:���.��)�~*�£�����ӎm��<�}�|��oTɈ�"����3G��3�J� ��`��q�6���o���%��p#W i
CrEI4���6E�:��$�1N�]mo����{�,�WF㥿���h�e�	k�ڳ�(���QT�:F�.�szh�3'#��ī�� �mC�p���QC`����,��bR�%��Q:� �X�Nu�pW��F�Yh��z\�e���h�1#�_�a����ε?��Ns�빂�G�MݦM2ܺ�$C0���$�3���Dp^9\aE�y�&3&ّa Ý�[��Ϩw����*�0S9j��_OT��B�(.Rd?O�1c=��iwϕ��o��\JG����|ϲ�ߧ���)?jo����M�6!���2���W�/���ѳ�&0�1 ���x=�@Ή r��}5�b
�6�u+hüh��n,Z����uscq��_�F�~'�d�l}�X07�E���kDAc+W�������!���(�	��s �� �7���.-�ўH�r�&�0n�*�Qz׹frx�&�l��m���c��}�@�#�]�3`�f.p����6-b�07�Oo�r7w+7
:�WG�iX�EyOr1�x4eױTD=ez�b�k'Cuz��o��M��̬�_zɢ����ٕ'B�d��E)�%�e]�aO�C��C��C^����স�{p5����A|!����ݸ_,��rG@Y��V�t>�.�\��|��|>315և'q#v	9�T]�-�H�{��W�n�z~��rX�d,���������mF4�v�֊*�ʜ���V�	FF����-�7Y;�R*�&����;6f��&z�,�EqY�����7f��˾�8q	�O���콕Up� R�zϧ�s����2\^�V�E̡qw��ꩁ^ߦ�
�rW����g����E�f�c�QrNav�w�z��*g��ɧ�b����f��9�x��;���f�����q֋;�D�gO�m�h�V}3S}�ԹƤ*��r��Od��T{�Դ��?S�c,�2���*%�T
z/ՁT�&�oM1���B���P�H���� I�K`
2f*�Q#��TrY�X�����O���>Q�D��21��|!?7s��m��h��nbE��"���Jg������O���ͫ%��|JJ��}Jh��S�����v��"2'�C�4Ћ@��B�M��6B�V����iu����a\��������ˁP�o�4��M枹mL�G�����r�}���CN�e����-�ƾ-���%���嶚���`��}�p�C���M�v	���@&O0I���tEɑ��b�����s����c��@(����6��p��n�k��r^hL�"J�VL�	|�&��Fk5n���۞���[=��=�h!���x�,���d��2ifOP؃^���K��hX����T���P �Yŉ�)l(K7��*�Ȳ�A(��/L�&/�\xP���%1`�I���~:������A���KJ�9y҃$B����)�$ʈԬbA
+��?/�"���I�5��V����&�� ��f"R��>��,�lQ�!,�2-2Kv��ITjlt�ve��^����[QCoؗ���Ձ�3?�7�z�N��>������"�8�����M�q�!v�E�E�˖4������$ȁL+����>,�d��u��yٖf{���#!e<��& ј���_b�I^I!kQ��O��hWE��I>Ry��<�3:�[��^ӂ�1��2
4b�յwddd��M�FV�d�0&��ط+K2��8y��]II��ܻ��?�ٮ����ϑߔ�� �m\�;��|�b4י���|$鴦���Bm?�S�%>�����z��R�A��$�R۷�������U�G�G{�Zl��]Y���s��"$!�Dl���XZN¶��,�t(��jhjS����!�����o�=��`�%0Sh]"��/�(��Q�E<���:0�����V��C[���?Y�r��`�|����T��7�ye���<m'qj��bQ�˔���l0Z�{�u���3�m� �X�f{F+Җ�Cs���CPw=�ω5}l�~qݙl�WF�>��$�`��\=�Q�Y��t_�-�-(�m�'m�d{�.�L�9��Zk]?�[&R���f��uJ�6�ɠ��E(M��Q�F�-��zj1�U�L�b+hh��S�clAL��U](͞iЮ�Z������K��	ڹ�l~�]K��Cʱ��
2�2Eݦ�!��|��M����DDR)P�����rs���40�Z�|F���o!�.�PH%��(1J�	�$���%Y��=1Ih ���.<�M_f�ky�} V:ڂ
�or]�06z�����?�y.I�SAu0z����5���hZ� �hΧ�"j��� ��\�����{�A�Srlr�K@Mo�#��.
b\z�'<��x_�t\����3+Vx`p��]�BU�տ���l��S����'<d��Z_d4���^k\����V�r���>��r��w��� !{�W"<qu�\�׉=xw�~�r���i�8 ��W�8���+^ zϱ��j"�	���Yt��uB0T��z��L^p�v$Ґ�{a��\�87��a�bDd��K~�쇈:�n�]|NŠT&4(@�8�-'+��H$�TIYxաl�{y��$��	�������^��n�ȍ��b)�l�Z�a��s(��i�H��~54�-rڵ��h8�n�O��Pz�Ő.�j-P�@~?y����2��@H-U�5�k7i�����r<����R������B	�ߎ*N�����*ӓ�{TNS�Ό֋4=���Q2n%�a-kJ�p�F�h j�?=�1�f��Zmn(��g:iK��Z����h=�¤!mI�zv{l�c���UӁ�&�S욊�g��	�zL.���3{b���-`�D�x�q�w�(�L�z�	�g�<N�m���{j������dh�+O�����b�w�� �w�������i]ؗp�py1�8-�9�M'"W-���3y�A�)�cr��ߡ�g����aq��B#�A��Ӈ@��5O�N�}vO�����f���z��D�ѭd=�m���`Hp�An���X-ϙdK�3�$���/���(?F��`5��
�.&�
f]^��G�غ���ԡ�F�Z��eȺ�535��Á0�q�C3Dì�co*�E�.�-J)M�M��)����>11Yq�P���j���"aC*�m��9ٙ\�����8���%����.C��Mͪ�Ϭ.n(]���-L�OݳGj�7&�W.��O�ոRx4��).%�*�za��1����f���
Pw�Uz���������m�M�3�"��X���-E�
w���Ⲋ��o�2~[����5����~BD��H����� <�����
TA��Y��!�\c�-���:-Ņ-���k��!��	�,Q����,Y�'����)���ڒp��x�$:E9�_�ٜ�/&�P�E�6��������X�J"gE��iY5�5���&\�0JUi�)r��&�R�1�����58\��:f3 [9c���q&_���k�i�ֿ�;�������eiz,x���HH���/��iY;Oy:�:�^.HH$�_�/M��M$#���Q�ՉzO�2�m��/���د���R���p�K��P���F,e��]K��dQK�!�� ��׃�BP��U��X�"�u)ۏ-�~'�JM>��g6��uwV��N���?��x�a�?w�ζK lq�׊%��xT&A�eG�Y>�Ә�J,�����>W�o�C�*��Y\7��ӑC�_�0r���R2�m��`����k%>����p왺�L'o7�HR��iSj��7�̹����06|��rB�[��p�r��	��T����J����\ ZYɱ�0&�f\wT]LD�Xu�y��&J`%�/|�o�d�;Z���L)8$�C�[�L�fB���K˚�������9^�(>O<�}��uUQ4��ɲ�v��h=�Ӆ�/_>NE�x{�z���A�_Ȥ�'�u ���������.��氍�?������R�U�>I�Wm?�	�T!��{�,�%ކJI�R�iA��"k~�Ps���mi��c������L�J�l����Ă��An�V�^-^��c'�,���G
Zu�Z(�[8/��ḱJ�>��]2{0<@��l�{�WcA5��[�[�|F��A�\y,�p4�@ˣ��iYR� ��.�ݸ-[��/ڇw�Ƞs��}���C�դ>����nߙb���x�Ɔ��}����7gw`��Q�������C?)x���t&�!b�߰>�ڳ]�+��)��Z����������`!ɓ+������W��h��dt���l���0�z��c4/�X�X��Ti����lNrz�|�5j��.3�S7%�_����lp+7%G�#*"U�����~v��;�F�z��o��j��$Q/�x1�����~��b�d�yܶ��*[�YlR�T<n�ֽ�E��;��B݄c_H��*�ऍ�[5�2�Q�[M&�5O��[�~�/TV?WX�	��w6}�o�.��,�¦�&�_�����fձg�7|�>�Z�i:�T�}iN��E����;B�L�u��6���/�[/nC_�����$I���S�j�LF�W�L���Q�.�������&�� J��K���j�Oƶ��?P��2��%а�!�z��v1����?TV����ץؖ��EtP�����b���%���8�tǊ�~�l�A&��*�<�1��� ��M��.�2n]_�a(��o���gw�jaO1Ɓy�R�I'���@�l�騐i"�DC�"aGL{��:���o4�[%*���7M����*����t��Z�!B��Í�� ��0tӜ?�^+P�߶�f%�� ǣ���&;ݵ�K�/Yw|T�4>�2 (�߸��/N��t�c�_@�8�(g�0 ��,�X��q��G�:h��9B��f[���<�#����K��f����6d��%\�᝻2�n�{��+G~$u�~2���uFB;<7�����`�X��G��=9A��i��j���,�u�2�u��u!�`P�υ5��+F.Bs�3�N���Ɩ���p�'���˻���{|�見�Q�J��Md/>�PO�,�d\��ƽH��G߷r�jO�ȏq�D���l�%� �!i�?%5�:����{9�����.�O�0}9ٶ�tE�����@ �K/8x��<��q�|�]�:�	 �Z�m��$*ҨM,�s@����C'��4m���C�PjwЌ)F�%��Q��<�E�8�h���])�VR�9g�P�������C}B)_�.���^*�� 7$��vd���DB��*/m��S4/�d#�Hc,	�-_�ҏ@��є�lgftc���j]j(� �޾��B�kF�5E�\y�z���σ�6�4�:q�m�M֓'�Fk&=�|�-<���#�B!Y����{�W7�ݤ�Zy)�b��)~��6��]�Y���ox��mj �P�W��i�u��fr�rw���W>�?���_R�Iho���}˒�6l�>�;BĨ�6(�>�dE�A�8q=т���"�\"��%�x�ݭ�Jn���[��?�F�tQ��aϾ؉ĉ������M�~�xe.ޤԵE aOo߹
e����oNahL���P�n��`�nӕ�F�1����O~R�S���x�KZ03�`\�t�)�y7�����#�*H�?�|�yw^�Ap� yE��d��ӴI2Aaeg�B���2���l]�vM�\�L�����f@Ƀ���E]�0
�4mz9i�I�ycPՊɩ��ݖG�IdE���k�mW&4���.Gż"�	"EO�N���}T:���F��S��E�~x'9�f��I���e��2q�|��)^`!�\���7�fo|�����^x/7��M+�ͤ*������m&��R��� ��dfI��vt��?������΍�f���5��_��h����t!�A�?���<��a��/R��"�<0A���6M��(͈X�xS�e^��Yq˖�cN��6A1��U,�c��7���r:'|�i��a�i"@1 Vb8.���_�h�,��qw
���T������䭇tD�'�N��v�=x5��4�'�����Y����ٓBA��!��x �EU������Wכ���Z"�����\�<L�y���;^��:��cs���n�eVp�(k�,C��hC��LR �����/H�I|8j��F%_�Y�>_��H2����O���JQ�Ģ�uo���'9�u��X��*d�ӧ/Z����W�c����ύ�'ʺ���T��a����e|��d�ھ����9l"њ���vSl��)��e҆�|��K*�>��~w�0���B�(��ɣ���� �v;�l����;��p��ت�SsL� �
�ci�Kl����������]k��_E���;P�e�XD�����Q�mp��k����I�!%����)ss��>�aA���\<��e��:�w��l�O����e	&�����X���ы�nq�o���o�������tWX�r�bꊘ�t�&�9z��k���b�}x�բbJr<���'�r~n\v7�_*�"�l�Q`�䐬~:j?CQ�Qy�Y�
X٢H��N�Į��6;U�pJ��h��ȇ�K��-<<�q*�<1��y���X=��%F�g�J��o�d��ޭUu*<
�:�+9Jꀑ�6���4OLe�2���]*jټ���`>�8[
�SJ�(�O�,��'���A���i�Z������P��A�Qs�A��T�~p����q-s�� �,�#�&��fcK��C��b�G)O�״Gi :�X-�hYt\c�a���Q �����W������ ��L�KDk�ഈG�>]��� O����k1_{�cضKF��9B� G$1�.�҃�]��Y�0�ӤO�w!�3��Z�&�?�;��Pr����٪��=�1���x3�WW�E�����v��k58�{7��d��Zc�8vE�_��1bZ��ʉ�rĽ�&s{G��NT�DmDa��eϩ�4R�Op��
CD�a�#1����$ߪp<��茋�t(����L���J۾0w�/�͘�����-T����S�\�2�c|f�f���z���s)�~����xY�ey��Iɾ(�V��-�iǋ��?5~�E3��U��q�Z���-a\�͐��j��B�9�+��5|�����5�
��hJp<חh���@��㡆�<0ֳ���͝i.�:�������M+O�`Q���#���� >)Ś)����;w[�#�\ �j�e����K#E�����s1u�4��r*��U p������G��O��㳿�v�θE�B���$�v�AǦ���5o�&�ohw�˒�*Ry�*<Pv�g�p��j�����΄��������%4���Bՙ`Ⰽ5$����"±�@Ee\���t��je2A�C��p��,p��t�f�?>%y�ϧ��כf�l�♮")�[�@�Kn.�M�
��Nu�W��W�4t�Я�E���;$nݛXI�0pWx*���܊ׅ���W����S��U;� @U���&�z%�I<|�ʽ`��,�TV���`)-)ᯱ�fU!!pj�g/�#����$qў�88FS���ʶT�[��/��<q7Yz�U	���N��`#:޻���}�Y{��.�1ۓ�D&w�@�L�#)��TWG4*c��4G�{S7p�'k$��0&�7S��f���u-��ݾ�my����U��z�s�I��t
�Ce9���)Z��C�%��p�#�Ԏz{L�� �a�Q�I׺6c	6�y>u�vF6��n�6�� |??Id��jDCM���%D&�Т�Z��Ds�F��z�S��o���F�T�3ɖS������Y&[s��ӏ�-���K���U�%S���O��x� ��j�?V�h��G��Y-S�����l�s=�f�ā|��ct?�K�����n��Ź̾rS<�̱O�O��?�(w�D�o��B"�ե�P��b$�n\1מ:a�I�QL��� �]���%�U
�65b�ʩ��1x
&�������[�����0V9�g��\5�0[}J���D&�\}D<�_����pءǶ��2u,�����N�-Hv������nΨ�ʌu����Tg[�*j$80z!�^~���Gl����n��<�M;dG�^�ܝ;}]��wz�!h&al�e@�O�G�eLgTS������4n\��S�nE;UG�����T����N�#q���=��4�U'cPn$���t�2t��%�oʏ�iA��E�:�l��NzAi/#����}��
���p�I������y{��� _�y!3������}��}�H<N(�z/Y�Zr�L@-�}��s5�����k��J��4�֦���q�VW�M<̡���`�_SN��u�T�"o��;��Q��*�/����()���y6^nw�R�@HgR�B��䂯	)�:|s���V,��5p_��?e���`��7�w�P�f����,'�E,rz<��|&(���,p����%��N��ˉ��/j�P����=B�G+w�
�bE� �"k-�#	Y8�p��<�l�J�q��L�@C8$���{h1`�k�WGc|����Rm1'n�6a2��NI�m��T㽙�"RK���Y��I�K[�/�1q̽N�{��"b���Y �T�����@�}�Z!�X�QR;L�b4�5[JW��f�M\M)�4��i��w���y�띜~�w<��Ȥzߩ�tаOt)n6��*�O��6��_І�i��T�~��H��^k�J��~G&tFD�)J��{�4�� �$�y�`���9���B��a�2�0^L��."M̋}aK�#���MO&�J+qQ�2\ �4t����4�9����O�9���<2%y�|��Ӥl�L�w�E�2�:/칈����{��t��f�b͸qo�0��Z����i��>�M��� ��%�-�r�[���E;����g�8#��#ۈ��|�Z�9j� ͂l-�?��-3z��Ώ��<ͷ�^_��[.qA��y��V�w�d���	!��-+L0@l���Ɗ�N��́��9��wQ�*�u���c�������' "v4�����T�s������gi���*ae�d���k$m���P3d�[�o��B��:3H��T0k�.�������t\4P+��v}ѹӇ&��&H�N��Q��g��Ҕ
�^g�d*bh��y����Դ�d������	@�pNYg��hฌ���K֊�C��!�o��j/
�Z_�u�r��2�.sk�.( Bn���>%h��+�Jk԰���S��6�P����e��;�h�J����n9L��kn�W3���pIݱp�k���O,����3�ϟH�檕oԛ}��P��F�lF��X^�3br��]�j}�X=m�c�f�aV'�����!�m���UĨ+�Ě{�}S�/���������|��.�����5G�P+�ٓ�����m1b��(�������&Õp6Ҽ����/��_Ob�ӯP���=�Ou*|��_{̛�"``nQ߷�.h��,�� �������x �cz�Z���,�3�Lb���@�~#h��s`Cu���(X5_}0��-��C�ʨ~�!���G����-(��QѴl�F`D���`Z��z�תP�#7X���}xP"�)-����o"³Tl4�z
�,ħ�4�._���#?��rP&� �%������u��o�βI�C�����bki�S��n���)F�x�y���٭��T��L=[!�N�(y~���Oi�(/�	���X:�~�?��]��e6��\@�*T\jg��&��jedbapu������)v�!��!�N����q�S|KSM&:b��u[p��~��8� -��z�������O`NP1����c���j��+fC������l��yl&w3[u\�A��YX�m�^4k�fqT��n
��9�.8 N�ښ�z�4�D�K~����4:���jP��Y�Y��D0X&&9����ߘ_ha���<�F��O�۰ֶ�}����#Ŏ�ŏ7�:����K�kI���R��@��N����)}���J�e�̽+<�lL��8�_�{�Ҫ��c���W9���#-z������?���2����g�����.qq�����&�M7�m)j� ��Ժ2����a|�&p%������ ��a��$ݛ!�ǳ\W
�:�(Dʁ��Ӆ�KI�
����F�9�F�y>��=�ZB�1���x�ɸH��3-�/��lJ�U�T��G�n���n���e�d��,��������qk�9�Y�j��H�>�@]�o�d��κs��SQ2�g�ixuŠl�	L%XGth;1�"��������Dx|\�C<�[Q~Z�I���'��!���U�P��?�b;ʫfҐ��t1\�&�CșTa����}�C� aACmk�ەg���o9��[�7O�O�JG0Y&@{׷NxC���P��2��'Qi�<�V$m�%��(R��۴cl�wt����a� ��Sj��5LM| |��ғ���?@���A�W�Җ�Dx���kW�ז*�o�ę2�K������A�V�����;���RK?g��B�nI2���y�F/��e�k�R���{\u`�Q�I�E5�NW�R[ia)a�cvͺ�L7�Ǟm_�$ǃ�n��Q��}8��s`U��
��D�ރ��j1r1�9�/�8ř��F�y�[)a�k�*�������Z�?V(|"[��w&�p:9%��UȺG<hIE{F�}
���9���.�Ew��ޭ�?G����Dڰ�Y��K�Q���/E2=J*�ZH��k�
�[;(jfBW�g2}��b�:.�p� g���(��OW$>u+ [�)���v����ΪM�o��q@�;�ށ��wo��S�z�ϥ9~���4��s����p�V��93e�w��k���`�p�����p�dk�%9�3ޭ�g�q���,�-c�?��-��4O"1�
Y�y�d]��D�����<��[�}�̪Vb=�i�As�����_~�X-�|�|�W�k*%�$jE/�^@�D ���9��$$�u e��A�T��4�$'�Hh	�P���[O�\ҭ�"��1�?Jl��P/�2�G���.��G�!fTGL� ��>�*Dc �F-�������ww*�\|���nm��N{ӖvH^�q[��^ ��������X���Z���$���*��X���0y�������>�9R���K��� A�1n�*�w̉�յ�4��4��&���y7�ܢI�M���<�}�E�FJhȨ�*x�5kUBC�˕�u��z���(�7����t�^>xo��i��}"#�\i\y]�A!�������<z�<8����ߟ7��؛u.��~��8���>X��j�5<��K��t��
���g�J��Z�W�hvڕ����au�	'���~O���itiM�)���H-��Y*����7|�>��D�]wԾz��ܓ	����,͘�V��u&�U]a��&����}[��v�W�̪&ؔ�0u�XNJ��cey�ix�_1Y�˜��40���AkG-��sb��G)������j�.j|���Z|�����o��Z�+�{f���\BUoC#��`���^+���4�W��l��v\�m<(�j_X��~� -yxVj3?t��FAX/���Nbu=D>��T�9�[���+�?r�W�l���q� �@e�F����ܠ�>�b1mfᅓ�'1�1)x���x���z�༿P�E���;Tbo���bL��3��²�/����Ύ�;��X��8˚ѭpÛD���P%���`��:�%��U���"�*�d`��%�0#T�+9G+W���F��Fu�E=��r��O�Kֈ�Y�_�Mi�ȫ���獨h��+����o��ľ6~wV���cԻ�&`ia ��+ ��rc\�~L��L���J���!��ӄ����t&�x�c�F�J�� ��Ƴ�7�r���7������r#�����Ʋ�4�wEu����N,��>f`�����{�s^�{	��V�ͣ�lR�0�����V�)���R-�P�9��wGW�5��a��4K��2�����E�L���B�]l�/��v���߅v�@b�j�֡�Ȳ���Q�X$��;��l�5������wFVE�W�[�B��7��4냔�&�����y���Yb�|��C�	���2��SM�4[o 3���RN򲣲Tt  �ư��h��&h��(W�����ڐ>�������ޔ=����bq��~�t?Ѽ�8ҁ���;n�� �� r�����5�'3�lWC��$�Y�N���X���3�؉l��Kx�"N	����;{o�tK�{���i_}$�[�Df V�u���"L��hւ����Y��HT�=���V��Ie�1G�S�W�����dC��>��p�C��R��x��.��>37��(�����[q�b��"�at&��7��QBS�g��U����O�9v���A"&%�[��6iD��B�]�j@���Jo�͑�o�_���)���^���*B���a>�Ns��P��e��0~P\�m�<��h����׋e`KB?�r�5 �o���
cXMUD�3��흲���_s�s4E~o����`{�ǡ���TrU�i=͋jNp��Kض�U������'�����L�G�������\�gs2�U��"� �
�/�˻μ0��jK�&Ag+�H�����>c��ش6��bö���g#c�����1���+Ⰱ��}�M�Q�]����:c	����	�1=o<4'�]�l����X�&�$�͑� W}����c9F�V�'�Q*�Ks�/u�YU{/�\l��;!��� 9���j�}ڣg>猷��~�]��ǅ�9�p�r�f�ĺ�ݱ���K#j(�#<x�3=YE/]G�|9�#Z�� {=�^�;�/��x�r��i�fn������I�~_�	%��M� �2��	�ߠv~�p�ʯMNSu���T��9^)��g�>�9�IK��)�zY^;W4z�~�,M�ؕ,+�'h�o�S�3�)�hg]�}9���ݦ#����y:KI|���s|�8�o�r�K_ �J�
�UO?E�5��L��W��m|+�o�M�1~��+�����,V:>��ĩT����@|�R�rL�*|�<Z<K�`��O�M����\�9CR[	��D��<�|�C�v>�\u�=)��Q��{ۻ��/r��n��m�K�#*r�È���i=��~{3�=�T����ef�Q������nS���j]u�YZ�p��M��h{�eg�J)��_�ڌ�X+�t6����[��ѫ�{x{�n��3��Ό�;��pD��0{����,�aTym=5B�ʆ^c�7�_��k��':�������&j�0X��!n�"\+��H����\O94�f.�X���҄oּ9T҃��K�M�nV�{=�����h�W�>Z���*&�F���Z�7o9�@v6�M�4im�I��	�d�9��j���u>M�,��ɖc�1A�Jvp���,���0cd��cn	�@Ը��`,;A��1l�+����(��GI����p&�΀���8u�~�E�߉h�����m�, @h���g�Ѻ�󸧜:�׈�"�D�j$gG��H�[7�(��E�j�ҏ�)>��r�X0���jp𜡒&�<�ǔȨ�\I������iF 8�
P3Ǐ���P�r��+�7�;���݄��3� �Hh�3z�38�璥��\w��&kv��?͉6��&�`��[i}M+�RE���C
�v�d���p-l����2��J�u��E�C���l�S�Z��K����v5]�����;bJB�����o�ǫ��!�a,��]�>⳦�a��j�d���B��g������q���E�,�-4҂p�z�:�O̲�lت#��� ��o���Կ�*_��˳�݈��i�e��h��F�3�>�t����S�]���3mxj'��5nb�b G%r��R��O��1�*)ە�
��/t����R�{v'4�o��S14�z ��e��,5���f��3)ۛ3���3�|��K���
��oF�n&ă�_k-<����.���D�ɾ}��(X^ZKpN�Әn����x����,fl�}�����xοeg/�<�0SI!��v��.�W_�;��c��
<�葩����(�)�V�=��.��f�^���w��@�3�Q+�������\����v�����t�-E4��JZ�7���B��(��:$:�r��RA}4�H�����c�ɔ\��.\�u4%7�%5��xt��,Zr�^IPi�O�F p��%�i�m��zm��V����ĥ*���@��|<q��K�r�ِ.$%B9�#0���4�4v8ۥJUō��ZJ���CO��::-����ፁ�[W	qN�~`�e3�Z��Cu�P�w��S�+�N�B(����!EԸ�d�Z�@y��x�� #�[8�>�0���u/E�W�b��d�k��p��μꫧ��Uw}q�uk��y�o�x�m`4�U�wD$�7�q؆�
���������I]7�������&��@�>R�U�:�ηC,�Gn0��uE�}P؅�a�A��*��� ��%_���V �<�A�i����&�3V���o�x�P��pvп�O�m�wz�/Z�P֔�=oZ��z��,��.
�=`Ŷ�9�/����d��_R���B��?�����)��:�-�8�漖]~`.3.B!�����<U�.�B#a	(��f� �;�-�����-�:��}T|#'7ˏ�U�F�
f$�6y�BQ&>�]����V�9�a�	;�֯M��'�$��w@�اw���h����-<tMt��OG8[J�IvG�JV�5��[f�P���hS����xw��;����<d�[��p��^��ź ����
�h��L%�>$��w�'`��G�	X|�^(�w��e�w�ׁR��<&��';�����P��1�����A�(.!�9m[���"	�|J-
H>[n��85���/��;-��Y�b}�������v�����V���k\������W�����(%�a�m���V��^�)��D{����	�����q9@�ߋ곎&�ݮ��?��5�S��\r]L��WX;�K/�?SID
"���-��,9|I��7L ��AnH�ZeI;4��ۖ�$O��I�.b�*��[�|
	]mh&��4�eN�$v��]{�Ѹƴ��_cc\S-�.��%~��הe�ð�L�V�hns`��c�Q��c���SBH!m����d�
;����H#�ʗ�.w07�@�����#"�x���o|Ӣ{��@b���h~
)ԟ��Xd��]���MV���'Mm�H��q��v4�꿣�'�������\��H^5�Q�M�1��Ř��f ��p;�6>�KĎ�l�.E���N��핍��Qm�j*�F`�3U*d�E9VqV���ʱ��|¹TS!�#��>�o��զ��*:Ǚ�Q7(iV|���h#���<Uh쩳���v����pc�P�B�8h��3�`��K�v��9R!��6�&X")�&��Y;\C��(��cb>��&�D� �7;:$��{�z�C�Q�u�l��YL�r��k��f(,Xq��}8t �>o
}��ҽ��Y�#l=�;�u�p�	�|C��^[��}�݈_�.�D�o*�
UQ�0Ƃ�|�+]�}��qè0�Y.��z���CL��tS�p���g�!i�ͪ���HC'&�}7F`���}OǊ���wR���H~S^�'�N�q^G:���Y�e8���D���O�T�<\���-\j2kZu������{�7+��*ߤ���FC���x���}1�,�1�r�bbܻ
"�z�V�E�\� ���̞RA$��Y4���Iˊ�	�}����M�m�����������!�w żd�66��_h)�)
�n���1�G�;e'�,\����O����<��iٯ- ���o#�ὼ�I%���m*Aݲ���`@^���X��@*���a	��5��*����#y<ﹷ'�G����+�?�O,�>�0z	�(�jg\��n�D*��}�Չq�[�R��K�R2��j:�����/h�PLh������s�Ib�6b��r L{�k�{d�zR9}��&̀�똕������1%Ҕ�c�0j-c	�T�|�P���S���0�etFl?���'�ZL%@��]S'�bbZj����O���� �A�Ѕ�j)(�#ؑ���݆R�o��Ppe�dM�S�F�8�E�0}�ne:;�b�egd�1@3�{�!U�a���T���i}�	�����|�˘���[J����V�W��&5�F��)����<��K1CƝ��
�|rZ.1�i�2�a�;�� �3�dW53hM��`*��|�����A�+j�]�y��޿Rz� ���K�����8�F�*9��-�*��|J���Jȶt�F#V��c�o8y����\�����tf煏j��=9S�~�h��k��Pl���o&{���B�Ͽ<'`��i0�\�����	�_s��}m����6FY&���wYq��[�L�\P�� |���x�6�ʃ���5�6�d�A�d�\A�3�.
�������G&rf��&&�nAn�k�o��0�S��ծ�{ڕ���т7����b+��Z��}���f�X�x�����͆Z��x���[�ylc��x\V�'Z�U^:0�����N�t��nJ4�eq��1k����P�cA*>W���d���v�Չfg�g"pO��f�\�	�k<��+��lH��S�.�R.;���syf��R(�Ff�,mn3ƕLA]��Qe�T�ȵ��8�8�F����di�u���h�q|���қ<@��LhF�5;�<u�kBw|�2q�n{���J�CȢ\\�.�L��y��,�Ď�_�˫�
���9��������˾�TT7��J۾�:O��S��n���N�P��s���([�k�D���ӑ	�#��w�d�ؖ���q��f�d���I���"L�
I޵P�`��:���*m�ES���lTL#��˴��V=5뷙�'���k�~��Lo�LJa�r	,�_Dc��Kj��lT]K!$�)K��CA�*�QqvM%.���:F��AԟB����*�j9r�*�/�v�^75*��?��5y�KsV�Am��'a=�_@��]�8 �t�]a�\�Od�y�8���#��< 	�ɬx3K˜��ruj\_��$��&�9�\�`��i����-��Fz�~gмfB�$$V��k�v�.:	���Tn-5��S�,��:���z�x�v�{5�p`��F���=��^��ŧQ�O����ugmaD^)�Z���UN�S6|z&R���7������R� �#�+�{9��#r���(j��¶/��b��u�.d�O3)��9����y�a�O��R�D���*Wc�1�I#�xM�l3U���t>���e`\�(v8<{�р
�p�T��=	`����#Tu����Sub U��UCԪL���A����@w��{�����!��W����{(柍��a�>WaQ��Z{��l�l��,�;z��,P@�U�欄����h�C��i��J���C�m��lq�D���Ps���Dw�x�è�9�8 o�'J��	�zV��]j�%"�^k�P��-�Ž�z��l�|�D�c�˵Ъ��gr^�G~F~�8O��d��_�g<K��-�7 z[Ҁ�e�xG������X8���P��_)T���RP�:.��5�r�.��h�V������P�x�w}oD�K�@�:��@!^X�dS�6���d][�&�V�C�s���;Qi̎�^�ER�Њ�ym��幬���=�a@�6}�
p�~�D��5���ܚ��)(X� ��vI�6~�P�v,	}��jYYvO>���Y�̗�,�:7��ʡ��=�'���m�+u�q��{?]�?�����os�a�ŝ�PuY�:��QB�n5�(�ds��;Yv�(>����Bk)�m�5��4X��H��&���;��u�3����#Z-�=�4��u����O3��{kg���@�6�k��o�~�"E��)�
�)+I�4[�5�?>Ie��?���޾k����*+Z��zVf���d���u﷝��4:�<��#����\:�4��n��#�GZ\j���pv����#��[�ě&��z*�w�j��O�}�~x^��o��Z�-�8���V����W����������q(#�;�_�T�
9l�������2s��Q�1󖴾�kKO��z��ø�.�Q(>t��f�&��߭Ah�u|�?�FM������p�j���c%ko?u�
A1h�]�7�@�9ѱ^zlҸ7���ɰ�qw��c�<�Z�'Ep�#kR�c�٥�}�D���Id�D�:����'�S۞���z�K����*(3�*QU�		�Y��ί��\�S�ut$������LDBu����:� �]z�C��8�7G"�� zH�����jJ%��O�|�2[���KE��A=�q�c�{I���K0����r�Ԥ��U�%�7��(v���v��	.д8Nbi�� ��z}e�ʞ�, �lnFa��MA����������{��7���D�h�<#���St��*a�E��/�.y�۰��a�{����]��=����Xէ?	���� ���,������=2V�nJz\���6�Hq����:�KT��{��V$.�擱�9��=�/.�! �Az�Y�Ŷ�1�`���aGVier��@P:iW�/��@ʥˣc	-Az0է�G����� �X��h�O-}O��6�aX�Ҩ��}B��} Vw�)*�3d��/�j�5��.2m�^sJK�c��s��������hK�
��	E뫗�0�K�:B�wD �]�.�T�ɞ�RԬ��1������ݩx�0�������y���Ȍ���Ō7F�<{f��mf��B]�`���Bg��z]-H4+K`�R�:��v<6	V��A/���<R�4e\��<%�z&�vf���s�\j�@�,ǉ��s���dsf{�KY��0#z��������?��̄�!� ,3̮�ߜ���NWR�Vpp�G�_�^�꒎8�vJ��d~�ER~(� q����l�Z�;�7�g�S��h�1!�z�J�~8���ίՏ8���{������Qs@�5g>��Kt5yG3�Y�r��:~�c��/u��[z����=H�n�ESV�h�z��d�i_`JT�QZ�����&����rz��6VI5��R�DJ��`K�sJ�*^��G��xf-�PcSh��{�ffǯS^R��z�NB�T��~�^'*���wO��t�����{ka�H���!|��9#��xJ��å�(kNz,;n�ԝ!~���lG'jϗf�6���\�E� ��^8i$��6ܛK��}�A#e��`���	F��g�������W�4"q\�;�㎣<'(��/�$o|OEF�BG�c!�,"�hL��~���,�w�bn$�wI��ko�J�d��Dյ�<\��x�U"�b����w�6\��\�
#��l�rE����рPȚR��ݧ9���2�ə�ٹ���J�gⵂ֔aEl4���9��J�Yy�:��uR��Ą�����2�nn�
��#�I���<�P�ם"�ڳKN�ʳ�´Y�h:X	��2�"y����wAfz�B�0;��I�ѣ�� �6���EG��]�P��*m�V�[�6�I�=^�"�l�j����g 'V�4k����E`N�a�B+f�a3��.��dm��d�D7��t!d����pi��a��^?��g�j侠��0'�w0b?R��h�z�¿<�ڃW�E����cC4'<h��H��Hu���-�'1V���ä����jY�Pkb?FdU8Z�ta~��w��
;M}�a�{�8Ҝ����M�&Z�p��|�n\Ǥ���;dWxxN�K֗�a�j�2�s;�*x1E)���-ְ�K���@�A��!D��ϭs���F�HH?;&�3/f�犡�P�Z��:��hG�>�g�4��X��=�����익���R�K�7��6�4��ä��Α�/Lr��ek��;E��y�|���A�S�n)�A�l�J�|PC�E����8"i{t ��#*T]���\3 �V��C�a(b)>������}m����tԶ���eϨ
��_��#et����q�_�t'���Wմ�.�C�Qa�SR�)��D��pr�A~�R=r���.r��VX%�&�ZOP�K�L�;w䶢6ֆ�*��in��d��{������6�y**�$X�wY�L$�!{��l�P��� �*j:���OMK�y�d�����ݸ]�wD2�=r��[����j�+�Ku�V� ���ο>�S��T-d֪
Bʊ�B��z/�o��;��GM�v��T�T����O������e/�O�ϥ����X�2�W��'����KӮ4 ]�,D'� �l�[��+=П:b��G��An�bG�IZ|��V���SĽ�"���'~�v2\��v	�a��.M1��t-�V�d�D�=H��⍞�LG{C�򐄔������|_�;��T��D6��,C�*4Ҿ��]��<��nQt6���&��N��~s������-��"��H�4�6%ۄ9��"{����3m�R�1j'W��L~]Y)i{�o�����]�g0��H��'�r��
�fj��X��PL�_�6Og�)1�Ydė�=e��C�\�dV���Ϗ��M:�r@9mxE�s�����?j���ы�a�s.�"��B<��������Jo�{��*�% xR�]�b�68
0�fNp���(�=h��mu��Z� 	��� �W��!��\� ��1��}��NE��P�!�b��4�N������pʉ���-��YcX٦Aaj�t�� vpK����\\�u++�]n�j��Sŷ���ð���
/V���M��~ȁ*1]I��4���O)�@ˎ�Zg����O�k����"�m���׍���X��<�~���c��U/����b3�
)ʉD�$���h1�D�u�pz��Pg��Z�)4�K�����ѿ��uCȁY����"yR�i��"TM�����2a@"3b����`��/e��qwv&�Yu��t42��P.ϧ�S���<��:�$Sd���5녋����γ�?�&�gj\#T�?�=K�^K���i'�cS�۽N�=nN�#k�zMq�}� ����_:��+���(��d�пI�%�岻���3��*�8�H�G��{�ނ�4j�!��d>Iz�Ka[��JZ���Q�e*�J>�JW�U�HJc:a6��p?�'����������Q�J�E6��8�/'����2ޞ�"VƇ}V�P��̕�D��::�>���}z� �o�F8�D��B�	w�F��}��١�N&�u�Ҁ��˪���>sM%s
�m%m�2G���ԓ���?۾�Vk���33Ѓ���4L����/Y�!�s�z��Ƌ���[�2�zY��������}�@*R*��z�Q�f�����v�|�K���Q��V~��3(-�gxL-t���^��˕����nIG��_����g4��D(��Z.�|awO�3ཐmpA��Ў����4nE���ɫJ@���T���2*��IDLB�fKo8�d�u��d�11	�2l7\��p��{�(��Z�:Y�d�3�Q������:�f�/]�wt"�}N#Xę���
��=���޲�&*�*{�� CsN���.	`z����fJZ��t9\����%t\��J�#��2��o]�Z�M1�O�"��a*��h�_���5:�˛M_���6C�4��U����1X�{&1x�&ňN[hy�Jt�4�ל�jX�lma�b�'<t�KI�H�&����<���ϙ����!S�QVƕr:�f�f�H�t��>k`��O��Ic}d��
M���ڸ����Tֶ�h57v�c��a��c$�ۿB�����d�B��,�o�<>�J�ɒ��<B\r~.�=f�!�UM���]ҿ�S��!v��|�g��!aB#�Ϟڡ)͵12�Z��,�CM�re5ڒ/|bH��o�m5z����5�����$��Z�_y�oby��"�ԫ��h�ֲĸ��*���/��ષ�o[9
����H�@�����H;���XZi�"	h*ױ��(�PݓD���%3��$�|�dQ���A�q��P�$�R�eNc���>0�>�6T��0�b����!�GHwŖl�K�p�#������v*�X����%t�Z@�@�L䁗?Cp����yA������Gb6�,29i����q����.D��GTA!̄�1M�&Țs"��ґjw��k�C���PN�6��
�L��Q鹄�4.���eh���ȩ�E�Zl��X=��b	c���z�5��E�Jk��2_
���8.��m��q:��WM��<-�ƪd�=�@g_���s�eo��6��������O:1�����&�a?2�G��/u�9Q�N�O�!���sb��R�Tmՠ=�;-��-#�w�+��Ջo�wPb@�_���- ֡�����ѣAlr3��%M	���9�>�A2^� y0�N��KBA w#'�Y4���UO�ˢ��s  ,a7�[з�\dT�zW:�;W�ґ�]�[O��1r��#V�)���2R�S��x��F����>�xŧ������W>k���Ҏ�	�`�N��x��/� ��K��s�ՖQ��%5�kX�1��V�N��{;�̾Y��?�| %����p��t5��6�h.�z�N���6�O0���'Շ�K���]�!?�s���`�Q�7������9O�2eU渦�nh~���{�t��U��2FH��]�Ϣt�x@�8O�S��.E{�Ο�l��9�I��GɑgR�I�y�}�L�~�i�~U|+����8��o�������p�tƥ��[���lc�9�ũ�ef��r3	��"�ڔk�<jz�����#��S#������&�@�P}��5�p���W�ꬃ~��������D֠u]HH���e|�ʾsL(�%�ʼa⑖%<F���~��Z�jDtc��V#����/Sa���$�}T(S��FI7�0O���I����ꝱ�C��	��}��LL%.�3A�e�a �i�^؀�?����`�[���&HH@�/�j�붴ąS	�	||�����9(ݳ��SzEN�C�9�Q�J��+g��z�W$p)���p��u�Z�3Y�7���`vF&3��Y<ʻ��F��>�����qO[��㬏,�mI����/�9p��O;cM\ݔ� �@���r�y�K�<�ݺwY�"��+���ژ�c^�=�Mٛ�(iBHl�6������w����s�^<�T�}��R��w��b�Q�&���
v�<�
�<��a49�V���<�[d���n��B, ���Ek+��Ζ����n#Y)�7��D�(:��P$�pvqy�e;$!/zz=�� ŬF":��s�|�X�:
{Sc'enOf�:��N}�Q�N�l�P��?��YvC#�+�:,lQ��\�/'����Y@��F�`J�$`�M�|��ʠ�P4�L�ؕ�Ԫ���'sy�">���X���=9]>y{�8��rQ�*k�s>#�.�D���ĭk��X�z������¢�y_@���研Q��/�Pܸ�Qb��e�� Z����S��,Ź8n:I{+��E�o��?%���������@FI�W��ϫ��e�3vlɨqLt)ZX�QɼF�� ����+����̭�=��\��1�<���3�v?����p���yt��
	��ߟ$�-�kfD����S�Z!j�M��%�#<��w��:Md��#O�+�X�+� ��/�d}�\ @|���[';�@n.��=����˹(.��gw<޳�yT�sN����6�H�ih:�����pap���)�ba�=��/{V�������?Z�ձ8�",Og/�E(g�X9�����,؛j������3G9�̒KGՅ<���KpI�*|V�B�C�ܤn[Ě��H��k#�C�7���;y��-���dڏ3nk�v(�q��P��L4���P^3�fJ&f��SUב�/~~���J�����L�v�8l���y ��6Z�.��[5;ߗ��o3<���R�P�7����*h�F8gI�ײ z���=z ���>��Ӝ��=�(���Jttr���8�h��C(��IO���\il�Mg�3\Cu�f�Ht#���8NGLESW�R��p�i���	��冻��R
���tgvGE�ao%����!q��T��}}c7�r�����e�L��sݦW]PY�sh���^#�Qy���ũ�-�^�BK����Zk��L�e�\	��r��ݣ�@���Z�v�`Z1�4��u��1-v[{\#���Bd�x.r�	g��������I�>/�@Ԛ.�`w��h��Ȗi]���HB�.19�gc�w�fU�������1���iQk��$�����B\��W[�Y$c$���gx��U�6X�ُ�S��=A�H~��h��x[.Uk\j����&�!p�?�f�*6_��/�\�r�l�t8B��lx�99.�Xv�y�Ua�=��Tcr���L��@�]��Q�Q�8.�-1"ٰ���v�r��Ne�	ZS�&��JPS�^4��
�/��z������wp�	܆(o�x��3;�:a������%鵠xTi�����Gtm���T9�Yދ��9bW�û�-����߾#�t0�4%�����֚&��h�.��7� ���zJVb#��h�7�����0�=F���t{��ڣ�C����TU���v[U�		��8�֖d��Aɠ�G½Lk�$��2��=ҏFg5b�o��:�F�O>�y�ip��>~X�V5��mS���
�A?����nZ��D}
���L���}h����i�.rk\�[�7bJ"��o�շN��:p�Z��S�*[ ՠ����S�|'��[/����tf[�)f|��dEOt�^��P�~�	;]%�LW����@��V@"�������Ԣ�t�̊���	�Y,9I��6�+�bo��)P��wd�Ct��
�e�i��h��j��	ͳn�`Γ��悇��#ۼD妲�1�Wm���"�,����$�q$�(-x�^h�ӏp\
�%�ʭ���sO܁�]� 5����h�j�:��eKG�n�B0�C �j�3�3csh=�+z�\�T-++O�9�-����.��/X�kMC�`�~�m��`�h%a5׈˲�g(�ȹ�6�"-�x��eT��3�K��S\Y�%&Ah��}��$��{�
��Ι�� �����,�3�ԡ 1��������"�4{����B�ߒp#h"d|�6�@�b����r��/Ӿ��A.�3ܬ�e�mx����f���uMM�G7�9� ~�MzV!z���N��=� 2��)Nz�V�y��%uG�C��s�f7+��i��+v�^ݨ ��ܞ��%9W]���dB�r�PlE7c�^�Y>pc�P
��qs{�B�u�R(C*���z�z�^��Kb�H�C��:�j��\c�v�JT�h�!���XI����<9��ӎ��ڱ�K*����{�SfzZb�~�ZͶt�w[g����U�Z��#̦�A�)V����q��2�:��c�%x����m]��ߢ:�!{2�l/���b�A%�B�hمsl�k%��U�G����mf�P�"�c��<E�7��v`� @]3q�-���lD��ⶴ�)2��W����iAN���sMT�/�>n�7->~-�۹glR���o=���Q��9�z����.�׾�u��zS���3�]�1��ܭ��~��N)$���E,zҐ����±l�7���'1Mlu6��� �Mi�fڴ�oe�e%�9y"
]�Ƈr����;;�n)��XL�ȋ���=B��L�^�a���K!��a�$��Et"�^ň�͐W鸳���)�\y�����uE>�;'��� *�3Wc	l�����,HE,H�{�!q���I���٠#��������L��3Xe�V_O
��t�_!�=�����y.��?�z`�+�p���L��ţ�L!����>�V���G��ڙ�bA3x����Z�Eߒ�h�3����]i#�oS��ZY⥐���XH�=��U��Am�bh"�j��٦��3�J%G���LT*��$�E��͠԰4��uo9;S��%��.�����zM��-�O�/��q^R����m=�~�P���[���s�������A �бgڴ%�)�7a��JԨ��&%tƄ��~t@,�,�л͹�/𭴀IY�t�]���z"�r)f������"r���*��pʭ�}]GE��ٰ�$n\��ĭ�B�K�a�V�u^��ZO��*�<C�ڸ����:$��ޮ���f�d$X;����ӎB?)Q-؊6/�g�k����	o�eLKI�=TL27�� ',47aS�¤v��yٙG�-�j,@����:d���
�����}���d��$�:��?=���77�`�Qn��D�����e�/�:ɬj���tO7�$|�M]m0���mY��a�m%�P�pͿ���U*mƃ��l.nM<�t->�r�܆g�����������%���M��i�2������2<f���E���cBm�@15�!�&i��t� k�e6�ˌ/�.��'����fT4)�ؽ]� �Uj�3��7�P3pf�q-���/�"oh��f�U�|�� �"��}j ��G%B�(�~Rba�Rj|�+��ʌ3'�7p�ED�H�I�:(�_����r���=�xb��0+"���*�1U��v4)�x�`�<\v�,��q��q���ڠ��d��[�wc�!Y����-^&�J��Ǐ@�%�B~=�oFAn�a��{`�9���L�y?�ِ���E3���t���>��n��@���"S�;�Z(��l�X���O�Io�ܴ�*�R����KC����{�*v��V!r+�*���*�չ�����Ny�P꿫���r��<)9R��3߲�;mx����b�,� ���&�� K��OF�_�X�K�e��'�k�]�;���΄�>��G�*R�)�5wv�3 �N�vǲ2B��#P�����T �ҹ�� (ܕ�XP]�,i�����M�i���eCpER��Vt�(�*��(~���V�@*��Y�c�t	!tO��_O�E����Q��"�Tl~ �1%���ZSd��y�D���°\zQ��\���^�t�^5kC���8@x�>�� 5���z��T�nVO�H���#��ՠj4w_��_�g*�>�G���p+���j�L�(�t2�)ҥ?�r E�M-��	�h����Z����Q�Y`�m��o�Y�l�+�j�ڭg�U��'�2m���-�C�Z�+�-�.�W�%��?ػo\�������^�	��7�vI�Vd���F�	�w�a��(FY�׏4Y�;b��&l���6���zB�ñ9%�b�>��&�j�0oƿ��:�[0k���k�pX����e!��+�#x^�����P����e�N������9[Hr-�S�74/���Jy�mf9�����*|�*+[W!\��Q��%��:W��Ĺҟ�tN���X��t*�� �������|)b�������޺@_�׿�xI��˔c�><�o6�k��!�.o��cຌ[��`p�3f�[���	�rkk��v	�c9��p��d�_3���Ѝ��M��Lb�\Zy'�e�%�2%�_��϶�D*p[��(
�,�>��d::���/f�S��\��䭻���0:N:�;d�'0ˁs�3�/���I���G�ӿ�����{?����Q�˲�8#UmM5��k��� ��^��zNbY�Th-r���}4v]��K΢D�R4�EkXz�RΖ�)�?a>V��h�F�A��:f+�-�q9#�W�쩨�;e2�D�0_� ��ぜS�Y5�!�dB$�^*$N ���w^ւF^�������2ٛ���l9f�qك\@���0�̎�����<5E�	���Wojbt��6L�~��=�A7��IY���gl��ʝd)�� '�����fL.2
B��������d�jv�f����|����6��.┖ƛ���N�����Y ��=����-�vHSF�_�������Cǜ��[~�bw0��J��ߪm��yٯ�,��%��~%��Uo��������i�oUfX���w2`�Vm`2w�xLS��aH]p4��E�%����0�Էc�����]�ߧ=G�oȞ��s���]@(y����`
�X��ñ�0S֍o�_ZF�����0L�任�����\����?=�Nɳ5������W�
��C�Y�kv�.�b4ߖj*�J^aO���?�]l�s�e�8O�[W�oc~0�u��"v�=��y���l�I引{��w�@C��)�m�Y�.�dI��{�������+q�cO�������ƿ�k��w�{�ô�#���ν���kApXe��_X��qkDc{#A���u�kr=̩���>�5L�D�;y��C�������0�E.�|H��q8�����:���)��V|x}�\�c��h� *d䞱�.���
b"�R�ِ�jpҎ}�c�����W1u��c��.�DNɢ�A��\�|R�Eۂ�馑��_���J�ٜڗ����Ō��ˎ�"�e�����%�wnDV��1�RG����zW�qeA�������kՓ}�,W|��כD@5����|�o{�y^5�[�z�<����]ۿ��m���NX��������w��J�dtU���Fƻ�����<�(�U�a�ve=���2L#C����$��� Ny��9s3�O�Nˍ��Z^�/2�11g
���p�f��6Eh<U��ߎ}gNxKk�j�\���7����c��ҮI�jq��?k�㕼����Ԣ�:�I[�LmЅӎ�S�c-nٱ���v������bͺtC����xŒ�pY�׺��s��͞+Fn��~�vG��H(x.�
:51h�L�O�׸-@E��>E9;<L!�O��j'�`m"#����0B�<]�d����ʄ�lrӲ�Ő˭ _��� �y��+![(��W��� "yp�) ��4 �۲W	o�Z���$���F?h{�s���;Dp)7@I'�Q�]��^V��Ɵz�]�+g<����2p���q؝�m&@h.5�[��o����I�䥝��zp�S#�hf���Wf�8(,�����B��;û�,���|Zg�0��y��j�*6���&nw[b�gŇd�� ��n���«��JW���i	P2"�`����HЧHOv�hY�ĥ�KR��}F�Md�;�w�"~�}^F �s)p�<59���F�t������#y��5��$��w�^:gm�9�
r/��G�<<5 K-��8��u�=P>쳢q�k'/�9���� �B'k=�#Ԋ$'l�ա^|��+�O+��x���v,pTQIмtn�ؚ����K�44~;7�U��Y�윫��D�ӹ�����9����CQ���~��:U��ш�1��o-� �Z7���R)�#�&��Ȇ��=�r5[���m�]f���!�����@o�vԗ��lϭR)gIm�9YL�G��)���/V�e�6$x�n>��Y�:h;d#B�%��5U�E��cj�v>V(_�g�`�>��Pp�6Ԋ?���XGM��'X�9n��nɿJo&�9�|iE|��
�1k���I�0'��*�2m��(�uS��4�3^��׌0Ⱥ���ĆV���2�c��'ș]��%�������z��Y6np8�E{�+���<�( v��6�
��}�����
1��a�6�Q��}0��������l6-^s��]Q�{�R�s�MW�/1k!G�"�v�D5GU��N�A�d���t�k�n�n���C%-�\M����u�)^�>����!�yj���َ
��U\�󰻔��|��O*�K�����@���u�gT=_�������N�4䄭�Ƀ���8��J�(�Wj�ހ3䮨c؃x��x(7�uB��7�~?���l}�b�֞�Uh�O4�c��)��{�Z�i�_����������Qm��*wI^�F��Lw��V��w�y��C��?�kH>�G�r�r�ZH��J �חJMO}��<�:��b#&��W�6�I�;��h�<�?�&O�_	P�����ג>2���>ag�Ś�;��3�֖����{�o8DQ'��s��n$[Q����_]Qk���ϴG-��/1�nu�,۲Z��{5��bЬЅ7��J\="!�Ĥ����J�S�Ĳ�dȦ��]{�/�l�˩����tÇH�	ڸ ���N��������5}���F7w>\ϖ�H����f�{�<��p�a��Z'�>Mc�.����K�4	��B�,CBM�+z��fg�"��5{���W�C��5Q��ݪHb��Q;EzN�;~�p�.�sT��.�.gh��h��m�p�̃�p�m���QFj�����!B��F}p��mN�!���k+��SX]�/��ۋ7�jx��a^}����}�_�l���f`b�m���=O@��2T�q�;#<P��W/Ҙx��\=�P�ЈL�ǒ58ACU��
v:Ff�y�H�%�i_TCw �K�{���q)�t�q�����q���8�rmD@�0�16�3�1�35tiG���a��&�;��N\M�Hs����,7g�j?8_��I�*S}�٘�&--�����L��� O��W�Q�r��2L�%�w�O����PW��>�x�<L?����ّa�~��UGR	,qiB{7�GBR3Ϛ8u�Q[V��V�u��N�<C��������y�fA���V�0��V�8�b%����hRu:���[>���;ʾE3Ux��G�v\�V��i��|�5�5F�i*���vIݪI�R�ۃ���6V(~�k��������0
���ܻڏg�Q����{n��s��JI��x�9-q�8i�"
���}���b���B�>���a$7@ӧ�rw/U�h�w�m�^0��zmv��Cʫ�Q���~
�R6a&>�%{ �8����4j�9���	��K�3�-���+)u��w_DP��R���l��'��gVʹ4�۸���o���϶1�$���G8��H�`����nn�y�`���P�G�N܁����S�{�N[����y7��'bӉ�ޏ6U��?M�z����wi?b��}��3�8n�"�D�U������z��,�ܰ�&��x�<�WX���f�M��o����[.F��/��bsA�Z��e�fI;�$��ACFz��3���i��4wG6�؟����pE6���ѹ.+��y7b�I.w��(����<4x��NqXu��lF�C�pmIZ,L��!g�.Mvf!f	Wē��,�m��>����i̦���*LӠ������]�;.>�fC_~sB��xd�c:N�5�@/f�io|����E��)7��g���&l�g˂�#�$�N]<VR�S�o�y3gܿqֳr	��&��mi��i���, �ޥ?�9zzs��Q�-��d��u��|���B}�R���ac��1ݩ�_);4�x
j��Kf�{�C�ҁ��Bƞ����"�ZVHp>%�Sm|��l���W$f�(�$�u"ga������oO_
-<�c�X3���%����W���<A�M�_�k��� �\�9▶ܿ_]��_c�xVQ{x=Y
��2�r~��φ�
�z�=H
������+̜�.I���8�Rᔪ���m���`I�ഽ巳��"��Uĩҽ̿+)U_: [
΅^C�zLƄ^^���S�g8��JQM�O^�#���rà~�W�FȪ�_�>�e䜊C:[������,I�{!+}�<��9�I�3e耂Ƿp�����k��X��f�dH�۟�
��d����)M�L���(������r-\ -��~�B��˒��9֖FHV)%l�����w�f_tؓK7b�����ݻ�� �{���_93o�L�S�FD�D�zנ+��[�\r�Y�m ���RҼH�P���V���;��2m'���_ϥu�����CSj�_�g�(r��kbv�W������K!z�N�,�ҧ��hs{�7�+�s>�H7�1�ŵrZ�zh��J�6 ��;C*�n�O1���Fp�m�#�P��5N�C�I���s_�˜M*�z��VC��KI-E��8ZX9��k�KQ�ɦ_������qfɺvY�ų�>�"��ά+�i�	X�I1GiI��m6/�L<�8 �W�H�=��U�'�ϗ�;@ �]�C���Hf�*[4�Z
��!q�����=���P���g`%�x��Ev�S_?�R��$�i��ǒ�7�XSn;���$�m�e����_�[ݝ*��ZE��it���'��s�4C|Gk�z��X�F`(T@3o��爘&a7!4<:�n�i�R&ЪЧ�2ϰp��Pu�^Z�(���)��M�?�u��p��V4K���@�]
@B{%��Th{B�(���¼qI<ށ.�7䊦�����P�0��
��a�)� ����fƃP�,�h4��'�/��Q����XW����u2�-Y_�V*9��+S
�zT�zWhc�5LȖ��ًD� ������S�+�����1��	��(�n�:wR���a��$ �DQ��k�y"�<�b`;����O�|�ꎣd=dH�`7h���2��~�BL<r�?��E\�������wY���+n�ӄ���t�0�?<.��X:
B��f7ّ��ˇ��x�����NTY�整�~��rO �A�ѻ���{����ɪ>*��N5@�aw�H�wB!�`Η�����Ġ�J��)�� ���֏.��T&72��G�;;�}�Yqos4=Ҝ���3�^u]�#Lh�ey;E5��ﻬ`;LM�, �?�ה�������(��m��p)�nπ��/���O���YbR���-�ٗ4_����͠� ����K�3A�������T����j�]j�P�D�`	�yg��lJ\̀�E�wH`�'�FЅ�O���!��7r�+���7����h�ߖ��"Kt`���o�:���b�qZ�k`�scj����oM�V �%>��;܊u��ڋ��A��.���~�/����'_�,�Ƶ;j��F������`�W*���ե����*Vr���.��~�����8����Z���2�P��A�6D�����b�g�}����&��߲��ף�E��D���گ��c�����i� ��8�A�!<���?���I+1+��1�P��ld����~3x�%���pK!���OG�?K�X|��{Uv�/�g�7ѹ���9�ژE�����FIةL�L�t��:�Z7���RĚ���4V<�)	��-٭?��,��a��G 4;����\�_q�aZh��ɒý���)?5�f%�0�v:2�ݨh�)s�P����z1')�r3xf^���C]�����-�+Y�6�����/������F���#�1�1� �\�_y���|���׶z&O�̴ĝ�#��U:S���,��H���e(�k��scnZY��CG���o��@TQ�^mfW��ގ���u����A�뒸�po�T��"w@���9�SS����9G[7��Zc�ʞ�zQuv�\�>���v@y5�	�(����'`�*�;�=���0�E�sm���w�C;��@��u�*�F�AݱO~����xl���0��C��"E�N�h�������[-Qgk�h,���U�q�H�;��ҥߥ�6;E�ܸ�U&�]��d"'8?�eh��7�5����;� �o�[୑*�����x2�Pb��������l��6c�5���2H��ic����6�б��\�"-ƻ"�HK��DƉ���C� 
p��9���N(�����]|nY³��	�B?K��E1<"������/]���HݑR;/'���I��B�2�҇�1  'f�+B��7~ŝ�Gy!��Q.�[u7d枋E���3��� f(w_f�]���J7�+�p�i�,?�`�,�vfn�;o�9����S��d��$pC�;|�q�׸~�y���s��Y��^�x�,GKxx �]����8-�^v��]ڣ�O���t�b���8lJS��7��P-�Ϫ���!�Xj-'L�n�?��^�����/8�9��8�m���#ۚk���7�_!<9MB!�
_��^,Z���0}�LaC���2��>��!�͟!tH:q��ڍ}&Ӻ�:��F6� z� QB}1����N�,�g֠|=|4��Bo�hw��O�*Q�o�m�9fy.Hh��]E<~w@�[�
~*Ҟ�/�@v)���2ou�Ar�D���Q��ʭ~��[[������B���sS�MâW������-������L�孙[Sڜq�q��6E��ʚ��Q*�#�'|�B9\�a� �B�\c�L���k�$R�!�BK��SQG2T�d�3�n��U���g�֒��D����h�K,"m��74+ �2�)���J�����B��J\A��`a�~�u�Ţ��$���>7:��I䜳�h��M֜��LJ���n.4'��'�)Y��*��#��5i�l!� Be�0������piXd�m�)�x��ף�@�cֆ��`]_Q����̦���á3�r���o����o�M��������!�@J�Dh���R���������Ҏ)P� ��o�9��3 :i����6h������!�I.pJT�f���Q�Xm��9w�s. 6;,��r	����)�<P�]ޤϐ���y/'4���$���=�DwD���zA��'g������S:B"]�d��m������Cn�l�{>ic�%��
�;QC�Ў�h�V�"ѻ�ɡҿ" �es��l�V��#��X1�L���Ӊk7�����b���O@���Q]��'g<$C��{�A4�/>�&�*9�Vc�(���Gs��}�\�7F��@�er�1s2��Ex	��M�2s[��.��=Fgܤ�.<g޻"�R�?�>z˱�Z��ͱ�_�7�K���ҕ#V��)�v�=��4 ��{P¿�=���
>�D�����B	�K�(5�@�wSR����}_e��؅��~�K�BMɠ�~����>M
V� �~q��øA�I�(/_���_|i��Rߚv�b��LU��>Bi3�nyh�U�w����E_��7���.�qۍ������j�ד<���.G�l���4uZ��=�d�2F�R`&�|S�̤S��#N*��A�%)�Nqt(������� �e�L���"ߙU�Hd=Dv�`�PN�Ow����}Q~vY������^9o����nVz9�B��k���@]y�%�v�jm��r�S��^���.��t��E�K���H����w�7�s���f_ȃ�����W�uw�����(�$Ȇ+R'�Ut��ZS��6�ehTi�t����v�挊�r������Ǧ�
;f�	��7j>p�{��8��_��6{��θ�v�1�Y˧Ѳ����ڄX��}�����b1oLCuxcJZ�:�x���|͘C�Ƅܜ�M���㹠C2?�x���g��:�ʬ `��F��n6$��[-@���D�����6zA��=��<��������mWǔ��7��QM:�]������ 
O��|�{��Qn�(t�.岓$�N;�#��h�NP҃�Fv6Brx�{��1S���Ҟ�W��dM����Ԥ�����,��8�2x��	�h�>��Z�K/�>v ������W��a��aȐ�wx��pÅ�rގ��y}�!�$�p'�KknP��`wyS�>��ۿ�Zw-G�0��?��{�7�)������:YK��!`ߊ�%�^�PW��w���ъ�8@��<��*Q��YQ�J�W�`�,E��Vo1P�mI^��X>�6�����Ji�2�ڰ���#�zlzjo�Y��:�l��*s/J[��Ut5[��� ���0�!��\9��-��f�C���4��[����(�y%X�CT���B5"J��6c�i����=����֓���խ��i�[��O�ۚE�`*�����2˲��������[b��픅(�T.zP��a~��	r�t�O�h�-�&Dr3��tu13&	N{�n���Nc�a�	L����uܷ&%W(�rFʶ��Wd϶��j�2�>CV�2��[(�B����hp-Q�I���\�SU(22��Td_Q���>!�������	uكw��b���J[���yθ�2C�Uw��#H�G���V$ȿ���e/�X~����B��qS�Ƒ��fxݨ��,I� ?4�p�B��cS�jX�0֠������J0��`Y�S	P%zv��&�-�*vN�xqM ��{ݴ�/#��b�3
�h�ڙsC)���So�E��1'|CN̽��l-��`�ЖYخbP���E��*���9O��\)�"cfQ�d[������ ��� �M��y녆ۨ� ���Q���$�۴� l�J�N����/CP��ký!�Ժ6��'N�2��ƫz�t��k4�6F!�������NF�ݵ[~s���[5�o3������s��Rㇽ����H��`�g�Af���� 4��~�=���@���� c8���.���8���#8-��A=�� �d�R-́�X�����F�񁶑�������b:P�'�j�gE~����)龍��Vp��'0�ha"(7_r˹�v(��@>�����|z4^�����\�L�缾3�/���#+V��2f�c�Tӈ��º�D{<�nr�@��?��exK j-
�*����ia�v�7�Ze]���86@߰@���@]}_+�}���R���MVp��^�y���ME�C� �9]R|:����^3]�)���L30������U��[,�0�w��<����!�BQn
����_���e���2%KbķD��[{U��� 뎘��I�ϧ)�J-���f��d�z���\�	�R�)�Ojt�]UP赍x�
����9f`���M��䵗PR�-�7���c���$���P�F�+Á�j����/n����T��,]B���3V�~����mF!	Lxz�'*���V0�]?B�΋�$��������]A��NV`���1tD$+FK�#�r��]��Ň���g?!�&M�\�ۜ��uBơ�2t�]>��~-�,xGu�`Ą"ҥ%����%I}��xJ��e��Z*)�m�C�U~����$"b����m��`4۱��H�e���{m���DFԻ}���>�WB�I�����p��.o���|��ܱ#��ǣ�����w������n�@3-a��٢��TmMZ��$ ��΍�60�� %�EX:�6A�~����Nz��`� ]�o�T�S���T�� �¹�J�������ΰ�K��&蘶�r�BXp?U,A6,�:���¾DP�tX���w���t�;!_��&|�����Y����8�=s��z8ۅ�PNP;䚵@Hcr$� ͒_��xl]��}ˌ�>�������#�z��[ X.����1�>�#�ys���\O-$s��·W��s�_K��==�A����Z[�L7�|q�Ө�pd�w�ʟr�q�(ۨg�5|b��(}�mۉ��S���_P8>X6_89*�a7c��/(j�&��rO������J�{��`�+��Ĝ���-���Nn<�N�Q�A>�;�dr��\���M����W��_��'w�U��6@�����_zK���u��g�����j�F7���y��[�q��=�k����I=*��(+Y�p��7E�Zߣ/�6��sq�LOP��-qȆ=����3�U���ػ$L[n�]f�5�=�O�|\Nۥ[�iL{����\`[T���g�(��*�5��<-*�I�)d��Z��!�^6��IN�2�#�eYek���$A�)p���\��h�0���	�d��wܥ�W��]�UG���.��r�[R�3���'M0��NM����@�{��~{�I���JUᝪo$Z�f�B'*�D �9k���R��pc:�}�� �������l���	s�4�Wu�� �d���
	��GO1���G��тn0R�|w����7)A$�!��Ha�%�i��7�,��)GƝ�dH&W�E�OB�W��fS��9b��x���u� 盕1/�ӈ��������*�wy�[������n�^GP���h���1��R����\�ZO45�G�5tP�<�p��\�ؕ�N):+$��l��x�uW}}���%߽�t�|�6v��s��U\ܲ�X��,D["��0���Bc1c�h��$L�}i��9�%�P�#��Di��j�Xp���
���Y
�;u2�$�fC�er�Y�/ә&�+RTp�h�w�*[X��-:�1��FWc<1MlP��{h�Ko�'ܞ^����P�DY��H�o���/�����g<�Qu�� 1�K߹�yx}����c@�|5�<�r�1  �M<�2�������[ݚ ��Yo�ZKA������A�>���n�ߒ|�}�&`�7ǚ,��>��F��4XR�f�a�BNO���0g�� ��i����$-�i.�A�1�!E�[����$�	\��{�l<������R!���,eA��YT�6���I7'(�y0Ec{�HF�K S���S�5F���Դ"�ၔ��2|f�Ɠ_���d�ᆉ[7��%�ކ5=\r��c�X��^~�gl��c�eln�&f����^Q݌Gc�ո!tR#����{���_,ia�ȶj]{��~x�y��׈�	��/Ļ��5`&֔����`.�B����9���m�Y������U����l��Ю6�6�����碒_��G�6�Պ���#J��0@�ϡ���W��o��6�Q
S�ã�_fe��>�����w��R�g۝����y?X�4��>���&a���?Щ�Vu;�#HG���s���P CpѪ�M���zu\���$ .ػ0B�J�5�xfP� o�oW0o�_�w�jI^ki*f->�+�G�/R�7��������a#v��p���v��H?��U��.ET�1ň�_$x(�PQ�m���Kޏ��6x�=��$��U��ꬽͰ��G<Q �t����B�*8�*< @�������&��@��n��3,o�X���(OW���KL���¤J<�-I�D��g�,�B_?�o���=���y�D���V%�T�l�@=?���,�/h>��ڤ��O�S�p��yv~�
/zW�������q�[�Y�q��>E��9�y��w��͞#e{iO���=P�@<d�����N��r�cs ȥ���<����뎥�ҫ5r���/.����e�1�Ƴl�����(�IO/�;k���:��L���Q�i������X?Ը"�C��ß�E�^����tZ<K}�O�)9� �Y��HPSܑyL�����]���� jh�����pps��`0
�7��H�[���FjZ<cĄu���Vȭ~xDCZ&c9��n���oTІ���&��<V�a��li>�/d�Y+b<%
�SO�J�k+p�Ď��W�8{`FZ��=1m��;X2����
�p����7�����i�=N�m�"`|e�©8C��.���sҌ�� H�V��%�0°��f���r�c�w��U��`�h�G�u���]��]�6t�V7`��l���RJ��ڹT��S�.v�'_I�<W��u�j�����ӹ�z;
��:B�5��4/}��p9܀l$��.�6�{Dpϱm��@kZ.bu���zk}�������F�����D��������Mt�-�}NMr���>-HxV�Z��͏A�r�$īK}[I�	���aPȘ*�z{?�c�ݗ�4Z�c������9����YfO�Ԉ�^�Ӡ��:O���(�;�����Me��E���ۅ/z��`7S��m���*���.��(䄙��,g�̃�iP;�S�AF.�s���w[Rh�6r�����9����UEO�NP5�z� ��Q�K�~��i.l�`�@K@�}z�S�T[�����'y���X��!4���N�+sx�d"�˘oM��?��@��:��@�7�l
�XC
���b�S2Q �3���8C�j�q��1b	6�C堰z�B3�M=d�D=����CC���?��]��R@���d��\��$�e����P-���<w����7�S�F��^5�%�,����,u���O��l�[]���\|	�o����W۾mU^��a��.s�� f�%ۛ�z�ϼ� 4T���;sj�2��K ��`�4�j%��R"�da��~<�Z$��C^��0����"�?ˣ�&�~b��}�8��0�F;�uY˃��[t����IA���
�O��9�L#h�Ox&��R��Xɞ���{���=x��6k�}��ZD-o_�lvZ�i�8�@,�Յ6o���d�����J��	ؠ���8�4P�!jһ��PФ#ޗ��q:4�瀊�*+
�?u���eM�G��v+���0,����6�����G8b�su�ٍ_n8�g�B���1����gjp�똽x� �?�My�����'N S��/rD�J��#�!O)F�����?�;���}L�ߵ��e%_�p�\ �9V2�[K�Q�u3��Mk�n�� q���YQ�+��w��0�E�{���T����Yw�6��0�7U!S�@�]e�U�dᐊ��]�����L+�G���d9��H,������2fi�B�տCw�*�֫\~xW�_�jE���3��^�ɞ�@�D^��x*��]A	n���s�����Q��-�!j#��A�lj��%҄���cV'��� �ƶ��43i�f*T�z �yK��i��{D�ŉΜ�j�T�o���:
�;��ޯ:��>�׋E4ܠ�(��)�%o��+jn�D�d�#�f�54�t�d�[����$�|�❺�F��w�Ĵ̣����1Kiq�Hz���'Io!�^b
M��#l�+��L��Ԩ���p��Wz����;8�Qb�D)�� �:/)"	O��_l��=��6TOԁ�öa]� ?�aG��T~
�S�#9�U1i�2-K
h,��3v`�o��� qcw` ��:K~o\�KW8u0s������X�V��8��	P���֗���v/������n�3rG��G�¦�U����'|�W�-�L{��$A�9��/��a'{h	�/��x�18!2�^����
��Q�JKC$�U�D=B+�� �0W�b�L�TU}���.�{�i%����uJ�z�'����gA�7��o�uȔ�{'i�d�_�brшE�!TL2���e�gy��w Da1�,�|� ��<�W=�'�7d� �1g-kOS��u4ZD="���6ٶ�~�����:���
�~cq�%����8CD���J>�=JU(!~Ee����6�{�#$ł/�uiv��1�$_45.�!;��-^y�iYз��U������=��1
���I$�C������E��t	��-\�"��e�B�e8�:�6ǏfS�ir�^�W��?�dej��;��!�uƑk-���v{��)~�~/��&4�� �5���i`�7�rC3Q ���Y�H��0�(�U����k<b�x��Tx�4�Գx�:���I��>��ש�?��T����nT��,@�7I�����d�rDzO�猂Y��`���zND���v����.�K��Ƙx>5��in%��tM���#C	��Bj��VqV=tݯ�D÷{�?툘��:��T!xs��1�%�0j���GB)Q�NdV�Ul�'B�M�QE�C7���_�ՃA?��|�B�uH�����1RFj�;�ߏ���%��D&����t�����"OI��h�Ò��Ҏ���sx����T�b�$.����T��#��M9H��v��E/�(e$Y?���|�o&�L С:�( ׂ�c��2�qo��������Sl��2����f�p���2s�F�r붿�����:�Wɢf��6S�I����b5h-�k���O�������Ȋ��D�G[���!�!��7i�n*��R���6�J�$4\=�Kd��&��#'�|�t�vۉy����F��7�j��G��@Ei��� �����$ǂig�2D��@Z��!�B��f���q���m��)��@>�d9�N���g����e�F2��ܧ�Wۚ�n�!����W��Z�S���B�k7��u��7Ο8*?X�xo�"$\VS�S�{�K�r��t�EQ�&bj������&T=�A������I�ݔ��gzAM��.^D'Im�λ�Q�=ڲ�_�h�e=`H�Y��5���� �>)Fe-7t���n\"�Y�˩��+G�*�gA�wYuRI?����-a��^���n��
v��&�h*߉��P�v0A黅q"��t�.�t�&��/F d�+�c��U�c|���]j�X9�z1���j�
,�:j�����X�%�!�cU�ۂ��̒��]�2���	��Z��J�vm&����]���w'x#W��M��|����%ay�����=���/��ٚK��	W�Y�,���*o���Q��o�!�����k�(Ӊ��aPFH�z���>�������YR��,\�c�������y����96k�Ut�n�焄���G��hJY�$��1�1�����r ͟��%���#ȋ�E�{�f�m�\�;6��W�~`�PO�M]�jҡ���K���VI`��Ɋk�=:��E�µ��Y��'4��<t$ f���+��i��G�A�X�C�"5�Pl����mѾ^�҃V�g���X��?�l� \_\7����	�4�)!e���*ӓ�"���z0&;C)��k����M��F�˪GQN�d)��9�x���$>�uA֔�zq	,��׋S�rU3���L?�% �����\��zX˻$��/ �y%y�!���l��PMfXW� �B��O���qn_��Յ:8�ކ��%a�6 u��FoT�ZʩR��-8�h�}��t�]�����>j��s�Y�4\�h\�E:ޔ��MFG�#
��<��k�D�X�'F����('���T�U�>n�b}uʿ�2��]���СU,R�g��j�뗬��:���-]��q��N-��՟����eQ��CmBt\u�٣�<"���[��B(/���%M�Y�2���jO�{�?PJ��9p��}"�1M�~[���<��-P�uU���0U�m�@0�O0�p��"���rxa��>C4�k�(�#t�?������!u�M"���vm�S���2 ��M�`�Y A~�T��G]J�`��ʪJ��<,w;�'B�m��)
�Qa[���dw������8������Ρno8�g�~3�\�X��Њ�1��R�Ԩ%u+���-�O+�{̭:�7~�xf^�cE�}��S�I�5,�%$&���ߴ>U��c�SMR-\�H�a�jZ v��K�]����[0H���_+�=��hjsO=1���#�ـ/a���!М��4���c�^��H���"F�R{ :!ncg5�
���,	�ߓCj鉇E�CBqJ}�	A�xH�k&�����$����me�n���_���D�]���yH�1TZ�����+�oaf��(q��-�͋M�H0M2�z�)��oIN�*���o������n�<�/s�>B�| ���5k4xD��I �$�ˀ��=N�����F�pm/M@�N�yR��BI�%5�O����ijI>���RѰ7�'���`��ߊ���> ���
M����s��}If�&݇*O�
(�����QnK���,ז
�pxoߚ�՗�-�?�}Xf��T�^�0���5-e���j?�$�I�ND�t�)� 	T�Kݑ.C��yw���qL�L��P���\l_�TА�����4��?�	�f@��łI*�z���]g�x��4� ݲ��9�����JȭC���u���k|���X���*��~�-Q��:��$肟$�b��iT��98����aj��_�s�6	�3�������
��C��7���f(�}ֆ��T��е>�/�yM��QR�4�! ����mݤ�����8�TKІ�@��1i{�,�!N���X&�U�q�6�>р�O���iuPY�
V���%Z�����E/˫"�˧控��8� R��S����w{�����u��6i8:���8+�c�ث�s;E�[��.w�)f���P;?����6'�p�7����!��9�+�)[5ʦ�6J��e��k�KD<s*�W@�U|�M��÷g�Cޏ6UF�N�i�� u{U���_Gx�����E��]j'`(��4g�ROK��帒�t{~��-������OŤe���Ss8r�4b��eA��bgk�r�3��D9�#UR��J'��� �c�jI�4�n���c�uk�p�Q��s�.0.cF>.9V�f:K�Q�����@41�� ��Rb��ׂ���R�>y�4a
�x�������Dv��+����G�Fi���:�	���4�'��5���B������6G�2=-x���dI���hx�U'Y�`�\j��87^�ҋ>��0��E%�)#��˘��v�S6�B��}N��ۿf����Ҁ�S�;�]X�K��YaJ�?e���(Cn��&�Grإ4�C����q'�7�G��[i��=���C�A����e�Z}���R6[��]�s����wc�@}��*���E�.�si����������1�@p����8F<�q0"�k����_�&�C�;�n�w��D1�\�&����ķ�qNf��2l�9!��B�@5�WKAH'�v��_)�eզ�;s⺬���)9G����2r������m�:�E@F��Ί5͂>���&���ZҰs�[Ԝ��$\Yd_UM�}�Ef���w�ΣTBZ��#��z�똌J:y��T7���:]�H_.���r�5�-�ou�җ�#���\
�d�w�<&��D�<�4�*Dq2r*t�o[� )���1w�3X�)rA�� P9HQtR}tk�\^�н�NI������$� �)P�@"��nD^�����k��y��jѿ�b�1�e�*�#�HTL�цQku��������8��k��D#�P
A��ob��'�
��bI���#�(�R�e�$�� [ �R� }�+C�*NӴ?~LO�]2�<�y�'f��K�f���J4MZ���$��W`�&�iw����V�P��D��y",JYV�����L�-�/;�������fj��?CZ(�u;4��{a֑v�.*><[&��;pQ2(g�����Q�aE�'��ًy(��⪳� W麛⯘(NQ�P��b�Bf��b�/?�r�!G�d-V�c�+&c|��}Ȼ��c03G�5b�#LBq}N̻D�O8�s�3}a�P�!���e��T����^�f��ͮ�=;g�0���L��}�1��������g �T����ͪiJ0��n��}���; �9�!�A���+%@�*?<�H�	ƒ��q)�z���/�-B����HN�R$�.�F0�����g��6G���W2�G%:���w��۱�M_�.���v�Yq��c�4~͢�&��Ε/Ҵ`_Hz��]��.�	��撃-juv���af[F,�茳�v�b���6@�������4u��QFǞ�W��+@'�-ޞ���pLF�ɨ���w]����Xٴ"@w�.>�fS��ǀOU��Iォ �#�H�����7M*��sڌ��Ũ��V,�a��
V�2��������e2�<�V��/jg�R� �/����C]<�o��7��ٝ���+_�&O��0����T̿#f|XY�/ʄ*|ގ'�ޠ�� �O�\�wR��b3%��k��x�0}������
�1���<�D��-�s�l����:��8��2��Ƽ�址�qr��-�2������o��ͭ��Ws�q�ԢO��j�� �y�Y�q�ʲ>�A�2@�C���%�flʣ�+>��iV��y�/��m���H���.2S���C�왕�po,wŃ�l4�V�Ù������sZM7��Z��z�{mk��ΫFHeW$R��`[i��4]�z}O<��"�E(�"6��\�3=�����O�ktomņ㉰4�Z��Y8Zm#Xzpv���SP��G[�{,��Ɯk����=o�����6��et��ُ�M�oϝ��|�ϭ-| +f'�FI"y[�b����G ��F�v������$�������T���pH�1KJ�*�pm*�w�L�t��wH��h�ݯC�dDHH2�X��c�]p��呙�+����.�q^Z�6ox�0�	
ο�9�<����O	2v���C����8~���a۹��W��"���V$Z��G��^�N:k;��ܣ�|�#�4w�tR���L&�v��f����/9�"��1ز�(A��$%�b��Q�P��y�Ȕ>�<e=�g�R��q⵶��\��z�W����ͤQ����Q��	�|�&��rXl��Dn���|���������>�`Je�(�Q+�z-�/�0G�1����Ͷ?���ûiۤ��"��| Z���Yf�|�M�-MB�0� e�VJC�}��<ٻl�������ڒSc޼��d�*2{6��ɬ����A?%-4/K�l�\Ll>���d��^�C��iս�p�2��3��6��Bc�$ײ���Jg�y���ݸj[�C���b��8�'���Ǳ�L=s��1��#��3#J1Q��*�w8����ZW��eq�XS��_��p rx#��44/n�3�ɒ�ݫ�c���!��!�ltn|��R���)�xw��qK,�+;�XYaG;��s�1a�һ��螜ԥ�7W@.K�����i���T�����}	�Gfןv-��HV�'�TnD�#���P˼��U��T#���`N��-� ���m�{�U�dW�%|6��]�?������_���aG�6�;��G��9)�E�AR�D���;Bi�*������K�U}���?�B�/��Lµ�4�x��/_o�$���g����:#$��N��A�E��qI�=���2ڀ{�(�X;�ʻ&z�$�͂����~��tk����W��y�1��0F׳��7�WJZQ��� ԉ°�\�+�5I�ZCR)pUq�|
�xe�o�I��N�B�������= �H8}˟��	��q��9�4�#���y,�"�c��@� �'.y��8����?-�.b���l�R񝕏��aW�����w{|�@X�Z�W����;�����b���-&��O���"Ь�E5X�5}�G�_�afI�ق�;�L��ڥh'r����U	�\;��J��:D*�9�	�\t����>K&:l��x��I�ø���b��͠�?@��U�.��y��`q/c�����~U.��5C��?��\��E:NYG�H��D�˘�5v����i�	��<���u[�N�,�/q�H�6 �	؎��Ά�l]�@�oI�AG�<L���=h��Br�}Z�3}�����9���j.o��Y��*<�x�X�7{|$6�f�M�mtEg�!Mf�0.�(��,H~*,!�ads����hX���������0����0�Y)��4� �1�w\d*�J�eB��˦�]�DQ�N�4�b�R0�[:n�`e��:t��Ҁz����bRR{�q�������v�r�N�����/ʭ��w��Nsrd����?�V�����,%��K��G1��������8i�?���~�JyG�m~�3�|�� 2�M*^�����;pH��Gp*�P�"r�7]7G':U`���ĹQ������a�u!kf渚o��8�Ȋ�S�0�LdE�6�ȭ6 -1:�{�n^Jv��]���\{T�s��Gk�s@{|�/��J�J�Io�Ţw�!�޷d����?�$d��?� ����@�y{�o? �ުut6K""���k�����	�֥_J�� $���:�׭�zn&V�d��������v�a.�|�G��u��;�"������8� ��j�u���x=�i�� �8��wۣV�ca�5N����~[J�
��}�fX��������{�5Н�xҦT�\���^g/0b��6T��Q�ȩ��fg,Dɷ�C>ߊ���@8���bu��wnďX�u��<��c��ϝ���-��p� ir���X��o�5"�)]�����&=�̗8���7�)L��<Vtm��0��b��:#L���$�qI�v�D��i�io4%���a�Q�����10@�?��T��R�X�"b3�\�d5,2n�)��~���Ar�<�e%�I�^#�O���9z�/ٍ�cё����-߅0�� ��^z:"2�V��!_���"c�WQk�Ҫ9a��(��"4"�$|�e�+	; ���pP@>R ���N\��<v1qח�X�����?�`���@�DD�WA��M��V������
��F,�i���`��1S�����X>��n� �Ӌ� �L�|䚣�6�Zbj;p@+P��ʧ]��%f>3�$u&�I;�Q�Θ��/��\n�$C�F=�\#�]�Ѡ-P���q0X�~��0�`���4� �jI��<��JIcY�I��9��A�)ZX5}�z<K)�L)>6CٺgA[�]��:ߙnj@��N֜F6֞`��2{%����!��p��^W�R����9�C�\\$�_X�6��X�f���P�����M��?�c�ۼ��?-�a�Z��J|�k�6TJP4��>��ß1��kis���BBWH�8D6�l�p�0�V����C�fu�r]�!���;�_-�#R3v�9g�1$��e��� �^�\��k�!s�<  ~"{��9h��.� �5]���}�h�e�a��wB2�������e��2%O{JcI:k.��jY���FS�?]���
D.�fyH�I~�[�AP\�C�&D�.�ߊv��+�2;�*<s�Y�������R��ɟxjyE�o+�:��ƌ�H��b6��Q���k�B�c�D+&����^ΗtZ&��!Y����k
3�C'N�G�[��ydx,�.i��SKԆS�d�0J�RxJ<�2la��g�Z񐰲M����*��a�?�j���&�煢9�y�&i���Q��H�
Bv�g�P拓��.��2W��p�ɳ4Օz�Iq�eOw�〷��Py����-�qNtO{z;�i�%tX�e�D3��!��CwDa����_��%����ݛl.Y�@�G�rP"N7���QtQ �7u�=���D�G�6L�kjL(�3^[_X�%�p�ހr(%��Tw�c��wDv����g��?ƀ��	%[�3�h3
�cć>�V�&����#�k"���'�>��81��<C��}Oh�Jʌ������8*T���w�X� "���pJ���A3����/2JFѻ��3tI��"��R�X���qJz�K,(e�x@�8���ު�(+0�"���#��7qޗ�QRL��Z�$�:�Kg�o�O�'0���6�����ɜn_���5[[z�׈!�v����qů��<�
1�@S����E���_$:��o���eV('{�l���B[c����p�z�+ںk3'�t˭Ŧ���#]j�D�+vl��t��,�xlj�3�����%�S��X�~`�`q����Q�jF
��_g�]�ऻЧDp�f��לeХ�W2��O����{�:�5��U���B²�,U|L C�_w�b՟_N��3�qG�M�\V:$�i�'FW�{6�?��НZ�ĕ��T�eeH�ٰ�dpYҐ����=W�!�����>�u=��=R�(BI�^�y6�D��
`x����h�D��t��k3j���FtG|��Hz��8(�t�YTT`�,�?#�R=7d$�ȡJRؗ,�I��4���ь`g���˽�E|��9-3�z��H��8��`Kg1�kX���~�J��-����t�GJM�a�e�~��R
��.� ,�[߭S��T��Ġ%�>�8��0[o����ն�E	.���۹8�1Z��U$��Ʀ��L'}ק��X�QI�v�"�f��l�����9V�}; �o��_G9�2O���4K�����.�*��m�g�Dz���w7پ�e۱O�>���x��_|����A�Ef;��j��d �!�L[�57n�S���I��DU��p�Ry���H�FsC�G�Ҽ����΋��7>\���g��5D���/a��,�:�H��n��KQ��K���@��A�a�F�odeR��}6*LE��*C��HO��+���]w��W���)��"H	�~S���P�R��IQ/m9�
��X�s ��k���Z_rB�i���,)�@WJ��U��?痶�<�]��F�Q#~�����g%����|���p�����
_>ۻ~�B��I'����+��Aқ>)'+��μ"<���
V^S�X��^ 2=.J0ٯ�PJ���af@!���m�a)9!ԁ~�qz�ӂ~䏒!�(�p��Y(���U4[�1 ړ�����=�$���8H��'��ִ2^ၙ~���s+:�3�]Q�8C<C���yx~�b����CB�mj/`��-������b'T��f5w�gE~FoP|����~$���Vڜ�U�)��͵V>�=ڹ��x�N�C�~XS�>#�e@@�AH�W��"��vU#��m�Y�`?�V@�����Z�Y�r�QA;���PK?��d�1�O�8���l/A�̆���ie���2u��L�b#sD�&R�ࡣˑi9�p�x��ˌs�\'[e�l�K�K.7˟�Ɓk�p����-n'd�K��у�~�f� |c I˙���n��--��ƙ��)�+��~�w�s�R|7��0��p����Kn�eK��w����b��@`��f�*�а{��%�w B`��I����M�8��p������>A���,��Ӊ��3I�����kw�BWu٧ө�����t�+�(�[Ź�j�%�G^i���3��9u-ڙk�Vt�zq6EIG�|�MFEhU�mB�R�ؚ}��e�8k����V��MEM1�سV��~�~�\���z"����&��G(� d���-=~T�\�Y��5D�5&~�t���&���;q.V�E\�w8Y��6<��G�Z!�ޒ�y\��p��)g:���Tk��[5"�[��.����&���|f�/�������ur�?W.-��i7����G����]�M|��K�vIV���_*^�)U�}�+3�#`�zS��8���-��#M�Q�R&߫���)jVE�~u<�{�׀��s,�A�n Akvwo/㟊oE��`�1��M��2z�7�ڋ81z0j�2�mƳ�ty�`+�Jg�H2��6������&�V"80��Ш�<�:�B��J�.�k�ܥtD#:���b�#�df[��"�赨rz=y~u�Ɨ��!0wK�~ti�~��ط3�v62}Z]���&qQ�/�K�1ҙ�R!�͎}'�F&�T�&U<��CR��(���U�8=pƪ;��Y3+�ET�~�W�6k/�J����C�9d����q�ѩT�h��ӝb{'���@���_���<�r8>s��� {��1�����zuޔ��Χ{���1l��;y:�3�h$��>0��T��6��<'�/���?D�z[`����\�ʌ�7�����qn���N���!��Q"�Pwн�?�[��4�ڣ�{w��۳���DR2<`�c��ڕ��	��~t��}�9�̆�Xr���+���W7�,�
5�C�a����bi��.s��*W�2�i��r��CS�m��`�&mTx춃�)#� ���=���̺Q_�4��ߔ�r���!�HP�s���Q�y	G�q�[Y�fn>��e�\�3ُJ}��_�5�����2b���i�#�?Fq��4U���D��&�s�Z ����O��3������7�P��0�;o�i����`Sp�I^��hR�ϙ��	g����\�b"�v
"���Y���l��������7����썅��]%�NV�_����>+s���hc�8O��q�}�����&S"�ݘv��sLI�ɗ-�v�\so�^c:���vϲu9��C��,�t:4�JҎ���n\̹�4E�����lk
=��������7�k�'���Es��~���9��;���ʘ�}(��MxW%�0�l�'�Y}�x�';�O{�C�2b��x�Ś���`�����x��Ih'�^�9/���m�UcCP!2��b�o ���̀��صu�#����_d(�L'�Y��ٳ,��j���\������{x��%���3p��ݞ�6�5k�XAȰ�q�v�䓞�����-�������uH�GWahmf�T�UL
��7�=K'�$�*�>��e3SJ1�j�$C@�煔z*��#��Q(�kA�����*��;������2p|#�Y/��Ћ l��cmur���jg*�0C�fn@��ߥ�G��c���2�8�	�O�$y�5[;�H4�\�?�*Ƙ}Ӻ��*s�i��X����$	\�Qa�F'��<9�l�Sz[���ߟu�_�<1x�}����S��!����p��0b���k����	��T^|%_���u��f�����'�Q˫��X����Bz�*�H�JD�H�~@�დs0d\��DT�
Ή�٨Kz+��S��� ��+V�����5���P�Bd��H��B��-.�k*�D~�u��4���y(v_�z����_�eF�MT����f�K����"`��é��Ǜ˦7�I²�L��;�Hܰ{�9<Q���u��g�7�D��n>�rR�w�w5�XY���G�Yo��v�U��4s9LJC��c�>�?N|����MaNDE��3�f�	�����gZ�פ9�H���W)��E舔�%����^̔&x��L#v���J��I�N��ϑ��+i�+�[I��~�Ѹ*�֮�wW����eރ%��V�e�D��90*xG�,��&�ܐT����k�������S*]�5��4��Շ\> ��D2��4�/���0�lf�R@ލ�WA�?A��6�y��ف���y�����.E�}2L���<@����㏙�U�3�]=���We,d���/9KO�q=F�C]�&�?���a��
�����a�R�|3�18�n�S-�O��aH�@�9S����T��{V4T�։�3�߸���ĝ.�Ԥ�q�,:O��kp8��@�� �c�wWQ���[O_��w���ސ�M{g6��y��YB������E'Q�<#w4f�� �߳�Uh��ߤbߴ�{�ӽ7�>�6�0�f�IW0z�؉�|!v�b;�	���5:H�Cn�x���]T`�d�kⴰ����
jE*��⫟ae��[;μޅ^�u�4��E<��)��q�(}A�����6�*��,�U-��I��`��8%�YL\�Z'g��s��a�8���#積�t�f��l�s��I钿��7w��8��N<��2�v���~��C��S�l�[U������}{��`�;�з�O<�R6�� EAT	Q���]�V�ʽ ���*�^�f_;�P~:���tS ��}'U��T	��	��r]-fɰ�U�oU܊�y�w�l7?��<��_���Х���uη�Hml���z��`�����Tݻ�H������@���y�
�4���HAמ4o��ί����T+��=��F�]+
���]o�I��a��)Z�w���û�g6��bL��8'��8�3��j�h���A=-�#�UtYFa�)����@a��$�*�+�kf�"孡�Xo�ʚ����x�1*�Q�@���R��9X0�w���k�i���Tf�����R�4E����ŅÓ���@�\����2	�S�!n[ٓs-��jB������$� �����g�s��K�:0�E�u��0���M��2�*���̛�ο.L��p�G#�V�Z�Q뙹o�57�Q=y1� Z�E
P�T&S�Z�����P?@\�GhK=��� 6�������30�ػ��x1��s�J/	<����V�¡uG�]�U�[�Cx�[Uc�&��:%�l��071�[��e6��'g0��u�pMBdZ:*A|yw��[$�Z����#Pj����j^������,��Q��;��}U°T����9#
&il1����������
��i��B�����;��;�TP��e�O���	�_yJ.T4J��d��zr�)��3$ѕ��{Mh���1���z��u���.s�L�A�qr��Ù�c��>�[�)<i�����$�	w�S�Nx����#�IN���Ƕ��*��]@7�{*�3��tD�l˱�1|G��O�_���yK�]2��:�$70��}�6i�+����|54���f���PG�-+�p�j�\��}륑�˘0��%�z&(S�c[�N��S媩�� ��ܛ��'��=��MP��~� ��S�� Y�j���������qU�:v���R~E��d��6.�Ϙ=)�29*U�-g����,{�����X���"�W�&E�mඏpb[��!���h/����� �ՠ�����^������t74Q�M\DnLG>�7�f���e�W���#��cf���u�&8i)Vuj�������-4&�!�k�;,u@I��#6N�1d�[Q�M��z%[|�g	I��˜��.(��*����m�hu<��mo��eIQ�ϩ��\}�+�nk�F�P��Y���:��ZB]<`����J��{L">�Q����Iv�7U9''e�{�+��T#*]3ni�o(�*Im9#��h� ��^�����"M�_��|hR�$��Ī=�B��Y\�;v��'̦ǶK����'���-D9��B�j4K�K�A=bk���Cj�.�ě������� !H.��/�L��lN��̆�~S���B������G�E���z3U�ߋPN�g�#�� ���4/Y�&�����D�?�	[��Ԫ�r13׶(	4�v{S�P0SR�|�9�����iI���Ead���ʒ;Zj�����*���<r ��e׸��gڢ�
�gO��{<�y%���,�����,hOL4�3���Z����3\\�B������n�vcM�e�~��"�����ްe)v���=5u�sY�^��-<E�1�{��֙�4�&�ی`���F��$�.�Pz�eI8dJa�Uz��/<{s���<�:R��W�£�՞_�믷F"�hI�Ac�~�`Oи��!bѺ1H]6DƂ�2��������e9�� ��U/�����ZX_Ew��v���:n+��0?���,�AГ�~�,e�'�M����c��7Rp��+��M��=1=�e_l؟�󖵡�]+��q��c��!�����m.)g)��\?�ۥ��3�� �����[V(��*!K5_�O���ڋ������NYy�")f;d,.P���5p�K ��Si� ��^ѯf��u0����w��"�V�?� �
�E�c㲩���W9
��o��-ͯZ1���F��d��:կivX�=Q(�'��������w�┌K� �£Ú@������n�(�(P�����2�-����F C�V�r߅�@Mg��s �y�������e6����sk}�y����A�#��yg�����=dl��b�Зy���c	� -M�'���K�N��҇#�
�0m�$:0-����w�b(+�I��b��9NZ�Th5Ƚa���ldv�9�t#�#?�js�R�\�A�ؾ�A( �����X:�Q���YM�d|34O/gd�d��XφR ��l<Gpd�F=���5���ZH��z��V������yD,�ڥн1��I4��=���Ʌi�~�h�y]ٖ���{���@^S����X9Ѽ��u�T����S�~�
jډ���}�g�,���1��ѽ��t��͎<Ǜe$�h��]�9�cK]k[��O(����*5��ˣ����Kh�������A���,I��ݘ��I�����EG��L��{IQ����{�]��G���H~��\ulO�=t�V�E�-*��~��N��ӡn����Ξe/�8���[��&�Gߤ�8:�|��ԧ7��U`�9����3��W�VT�W3��ow5�����d}&ۭ{L��?���}	H� ��� ��^"B�}j>U����r� {o�ֆ�Җ0!%jg0�Tt/��ѱ.i{4�T� ��#>I	Ǖ'ϖ�sK3�g�#/��C����qF1xa<��Z^t�Vᖺ���E�?����歼�n]|l�@#%�Y�k+��7���h��ۋ�-���7��_\l��'��'z��;�O>�犻xu*��S ��&�YB�Q>s5#�K֣��R�Bȵ��S
��!���pL6-[�_��<��#��F���A_X�
U����	���t��)��$�&F��LD���*�呷q��)=���.1�>S�ϐm� S:tG���3�	��[�z����nLb�C	c�
A�7�!�A>�U�޽.��Cu��76��Y�Nu����_������x�^{w�s=��;�,sя��x��D�<��ma5��.��)aI�CI/��������'w�cd,�f�'�����L2�0E��l�LJ3�D��x	b�"8�jH��ґ���w��7����Ϳ-=.��B��b�)�$�`cC0�sE��Lĺ���.�V��S-Q�h��ޯ�x��(��a�i4ѭ��7�T{̾�r����XM��['���B�5��+�'�.��w�!�	=�,�$s�[��:�k�mvy<.[t�;��pD�%W7��^��j���Ąa/��
#�@ۄ|���湢UӾ�9^3i������	!��y�:!�2���|���"0��ŵ��~!��<�`�|��N�S����J��`ҚRbn�A<
F�\r���N�"�%v��#g~e��1�G#��s�����	1j='���X����t6��n}%��syK�	��2Vϒ�ȧ �[��ȩ�߬���(w��n&pn��zH�`V���w����s�R]�l	�Dd�vG�W�%�\ݔ�̶v�©/�����Jo)L-AD.�L便��$[�a[����\ru�qF���{{QS�Yx���f�+��44K�T�9�4�4�ۡd�������K�V�i*�YA!�� z�|uѕ�T����@S�#1: s$�Y��;� v�?]o~7�nx�C��.lD�y�h?o@$!�oɉ�}��/h�܀6��x�>��Fx�H;
��U�{��e�n�v/)g�f�
�:��۟n6�4/-j�O	� ��i{��.��ϖ�Z�i|�qm���֌8�]�D�;١!{=�9��DĸY�Ew�k��$*�LD|?ã#~���̄��um�h0R�� ���-]Qэr���5dm���Z�������|�skH]�Z�_[D��''(��t����*��u�?�p��j���_>��2����4?�T�T귝��|�я���탭��W���t|]� 0KC��sp2#?#��-~�d���1EգsW��3�9���Q��0��j"�6Rl/�S|��i�;~��%�7&)��T wAeW�%fE���R]�)	{fV����k�v�%	U�I\!��p�Q]Ei��o�D�Z}�^Y��L(m�nu�yDw��LZ�8�s�:¢G"]�� ��z:<����ԑI�r��A�W�qw�1��+��d�Օ�����"�ʲ�����/���x�52��VL��b�5���(أA_O'�2�I:��yZ��ꁩ�t�`S��̎EW|�c�ac�CU��2��w���<s�xe�"�NM����ky`E�+߃��*�Ot)���2�_r�����y",<��~'D�g��<s�X$�Y4qeupl�����0���N.����ڂ�T�~�e�T)���.j�"�ĹO�%��']�|a�B��͏^q%�XikYC�h㰨VC�[�w_��#Y�o����X�DQ����>O�9�,qv?钚��C�͂D���V=��[�ڴ��Sy��Cܤ����6��Y�k�mSth
9S�:��P��B����BV;ߥ�F'��ewT~�K`�(��-�!M�4�h�Y�>��lV�l�C0G�ԑ�մ��;��$	��[�0h��uF�T�q��BK|�9��A�c�HY�I(�*��<��m���~�c��(�|��G�B!���/�S�s8�����!� �ՕFL��u�-����m1��d�)� 20�ǞԲX�����26M=6F�\V8_��4�2�H���������ovK̐ڝ�t9Ĭ�U�Kc&���QPB�#��U�->���P@��wH��v�j��FTN����w=�
�Ey>l&������n�~~�td~��۷!�Ҡ���2j"Q�����yY��Oy%9�^���v�?^v�d�m�F dM'�;���6�>�$ΟC��mr����Fqjeٳ�W�f��ɴs�i���e�Y-d"�l?�� v�G�M� 7t����*z�K������@is��,`N�rS��+uB,�67�7�cEN��d�1�U,��rث!������x�8^;W��߆����t5_��j0&40����b�N��Gc,.�\�|���]h��GZ���-^#��)&5l���)������EoF��[
p�k�j�:��������цYfT�x���?h��V�,�q����9ଜ��<"�y�4�'�`���Ÿx��H���C��D�,b$�>mw��eb������.�]�^A�7�$;
D���d��G!��l!KU���z�#5����Q����0t�!��� m���|��v,��	����s�� k���+�D~m;D�-;�I�66�gz
*o�B� ��&J�{	�����ҷE*� H��.H���8ک�CEc!A�+�nXI&N��M�dʍ߯_^ �H� ��æ�� �*C>�jg�bS�	Q��U�C�*���|��'Fa�������a
�j� �n=w��b�e�{X%�� ���x����<beK ���a���lGE��S�F d	��Aҟ����5#@�v-T�E�|��'��)���T�k��E�G������SRpZ��Iē5'��nQޑH荡��R=A8�&ʽ��Bs�zCQ�@4�Y��c4�.�oØ�u��Ŝ�#�5�Q��W�/�9sf��j�1S>8r��P��q�5��˚bzmk�����ɔ�Y[�� Sn�J#����QQ���Dma2�I��d@	S���0����."z�cE0�t�49�0G8�.�g�*�0������K����o]j]�����;E��@�Nȵ���d�Q<$�"�O�,�a�;ب�ԗ�)K�7N� ���ĊSB]4d�%�p��rKƦ<�wȚ�����9�WmBsG���]��a�q���8vIdF�\�`�Z��f��+����U�Q�g^\M��nmz�$���Tُ�"���}q�O�9*�Yn�B�������z�a[� �����:��3&x�	�� &d�ͷ����_p&��q�@Wd�KK���.�� HGuC��;]�<�_xMI4��y���|�<�E��5� ��*/�*S$p��D  *YƔ�Q��o?YV6g�$�9��"R�Ȳ�(�9�eޒ�|�S�ξ���T�.�`J_�sV�yX��2��p嶥����PmHB���R1;��B�k'�0_�c�b��G�}�����-TQU�QUF��7�W�՚��XW�Z]��d/���d�y9S�^Ʌw���\�8�]��ôc��E��s�U��t��c�p�Bvر��2]����=s����ۥ������[�Z �4�oˁ�@�B{w��wVh��0_�f��<�F�Z�^��T�d�[��.Q �"�n�dk�5�a��+���&�Ґ#�~��,��$.����^,��&����$�YNc=�h��\y�b��	cTM]u�=�"�4,f qg.�����F�dX�Ҩ���)3�4�7�3�28g�$���j�Rc�(��Ff�����f��J��#���-���c�Le�^v�lA�6@a��'��h�'E�}GJPX7&1 '���T}��n��6����s6��?2��|e�{�Wd��7ʚ�vh�6�IF5�0�_3�f���̦����i�!�c���A�L$�K|E� �Ġ�d��c'��C��k������>��x~?k��Y4���ΘYI�����f���y�a�����������8�@>DU��q�H�N]K�Ef�+�&7,ee�bI�o�î;s�k�/�SJ�]��r1����������ǚ�`��e��U�Y��$���W�F�㾸}�y��J���۾�RC��S�IR�=��'|w�G�
j���GT�T�&y6W�� Ï�M������%.��4�iLr/��Lò��U�/���D��/�Ns�Vj��Z���DTS_��l��s�384�����<Ȍ?.aW�si1����f3Px�6�pE��3ɮ�YEǳMi��~�oS��v���2�Ϻ��9���Ei�Qp�^���Kʘ����aB`P�/��@I��	i5�ɛ�7)�X����س�`I���US��$�O{VV����n����&�p�\0�I*���i��߇�r5�Cf$6�mR�s_�t��F����}���V�+��{\�����)�R�J�B��%�Q�f�Ӛ0w�-E¥|ƻh�]�/�.���PUh5��O@��<�w��^Us]h����A��^GM\Q����eUE�u,�qT�/��9�\��7�I�IM�ٌ��RJ$�.'hd��NI:������A Vޠ�S��`:n��D���g�M��7�Zܥ,c�G��-V�!�R�����ep�y��˃�0�"2%���|����>|&���J�]�2lG)lŕ.2g���m��DFz�܄��T�+	Y}�Z�P����D�/��ڞ�J��l	Ok$��a��Pܠ��k�T{"�(=��v������q���F��/z��4H=VԲ��$WW�ӠL"ȯ�����dK���������1�8�-��)��h~L�0�I�;.bF�c�/�솼�z#&6��N};eoeK���<���~�OS]�=@�z&�1h��q$"1����(-t���.���CUj�f�	�@+�NA)��7�����ĵ�
������A�y��|�8и��?�������$n2��5���?	z�f����*#�o��So� 0��ы0����~l�J��6���i����i�\@=P�5���{_p���!��S�/�^���}�'��ς`�����c�,."�%�)+B��n�nT
� �W�W��Bo�eے.��H4ZFv�4B"b�gH(�xR^2-��k��#&j��F&����m�~�'�9����&A�������s���ne��y[vb$j0��>d{պcޮ v�ߊE��Ͻ�AW{�4?�\�]��Cu�<
��u�ٓ��\�9:�\�6iUR�΅Pf��HC~M�U?2�.uS�#T��z�%����\��_Kl���RT�L|NHI��E����JaIt����x�2P�X�-�8�B�o d�y�3���0)�2����3q��nnsNFu_�����'pW���7�u�R/�;D�VMcOO{�$sUڣ�Vt�;�����Ni�Z�O
ɘz��@�ۃ��#�C�y��LRW��u���Ի#5g�Q���1=� )�B</΅}p�1v�%VQIƸ��8J�B9�0���Y�؈�� �]��r�K��B���f�
Mq���hCl�r��w�݉E!V��A.B�O<����B�o��ٍ��*�@^�pl�JFe�z@;����ZH�����F�QXt�,3񈸾ɹ������	�o��S )*��W�d&�J�^�'gGw�Ɯ3r���t�x���;RLB�ޜ#�gY%�^h��װe(�/���RZ���&"Ի)�uЉ�4-wb�?)&��k��+�ܭc؅�Ԛ^�S�l�w��*��k�rѵ%Ąߖ6����8'9.���ۂ��!�F-7�8��E�q�<�i��6��七-I9U�	EJO$�Br�c_׬ч���?��q�D_�1�n�G�'o�RZ���K �"HUݣ%Jt��|3:�;�8t��I�w�_r�O��=��O#V� 6/�c�q͹�9����([���	Hv�I=�iu�(�)�/��jT;BEe�x�.a >x��l�5�:+s1��.�w����b0,��a��ת�� �O\���EG�K�J �]O4@V������M�X�����[���R=uJ��֠�X�@�1.mU��� ��Z�'�^�%�Y���<��aP��S������3�8���j����7��=��-Q�,�Y���,�ڞ_�N����� ���N�A¥���4��ɔ�i�eǖv��6�4P����T�X�:Z�滑��Zܶ/x�9o���d+��!��+��1snךxEa���P�r7��Z�F�C~�g�j��vX)hcj?i ��R�A�����3�H��T�����I��S�M�Ƃ]�����c��	\92%�1�l����-B��I������BA$�r[;<U�.��̠=�d��,����:�L�.���� #��j e���]^o�#���?��5ݐr��
�F'c�K?�f�Ml�E�
)��8l�_��$xU!�8��sgE��h�Au��y�`F����Y�C���nd#,��hSo���x��h�׀hj_'��.T����{��	�/�lU��"������I�V	hO��(�	0�j#��@��6\U�S[��*��f\'4s`ޠݒ�p�ӏ�j���iG�[`a@at
�Z���Ȁ�h�8�`�^X)��:�{F9+�Ym $I-���4ff$s e|���4v�a���Y�h~{_�TDU���z@,�X�;	�:4�1������p+t�|���	m��.dIS%]���q�:�x�Qv�S+���Rs���$��y�<��#U�^ڷ0�e(�T��V�*��!�ae�������a o��t�Ӻ��-R�B��sF�r�>��1����A����3椰����8?$��ӥ,�R
;����/��>o��R�L���୿��cD`�+3c�'X�&�f!���ep_c�͛!��'���m^���<Q� ��l��@M�f����b$n��ϊ�P� O�$������K���0�#��>�Z��i�>9#��51!U��O��Q�m�9G�GL�Wn�Q-d�^z)�;?Q@�l;!�x�l�m����H��7���5V�O�YY�d<.�e�*�֓�7��"q�����u�#d��s��p!�qz#y>��6��n�\i�Y�0�ՐуN���Hz������Q8b�za�Irm������Д�vK��ֱD0��V�ɾ�Z;�Yr��7y��5O��W�bydTT񱈎ZGJ�X��nMv�Px���ч��OB3����wLՔ��S����^Z��i`ą~-Z=����S��K`��"�3�?)������R��6ĜU$�^�k=�<PY��ղ_΀eϖ�s:�,���ĵ�c�E)B��^��LZ||ѶIt���.�/Uȸ	l�s&������"�z�;~ErA�40��P�����e�����6c)�/Ș#1�����?ź�:ջ��!���C}0�"��r��;�Pl>��d�fbt$�N�\x|((�ggI-r#�-(7�җS7	�sL�;��.�X%XU5c�q7���Q�����u�����s턱�ږ��6�#g��!�����o�'�6�x��*�4�KT���<�����kXW1LԎ��ޕī�CN!��H�Dc��N����\E<������}����Kh1Z�#J%��1����rBx�@�d4e+Y�^�#�Tz�D���6���"��	V��!����G��=����E�F���C� �k�5aIڣ�C��S�g%)91��^��HA"�{hm`S������@��Sf�bo���LҚ��Y���}�����C@�^�$M�r��ʷ����E?��V�aKL#!��
Z����&�Hǉ����l��3��P�m�@���ՙ0*-5��J��wWʟ��t�mϺ���&�AIf���1L�A��ڐ������4�#��p�8�Ug��Pyj2�m,'�l����� V�^oO�9B�z˵�c�ڱ�9?�,@ZY�H���5
�6�I�N�XNE�֏��)�W�˛�m{�h�8�:�ǆ�1G���ӣ���+�����{8E_���Z`��?2���H�^��D3�kh��h@9*�r�8���62����p�Q�Ie�~q��K��$����	d�BBT���������QW^ދH�.�5ʘ��6�R����v��1����'b�O$�q�����s�G���g��Ȅ�Zퟮ�>��vxӒE�G���uڂ�h�z���26���T���R&�t�ctR����L�G W��W<n$ ~�f�S">cb��M{��X͡�D���K� �S�?���iB��<�k}:m�ᄬ�����}����u��=%|�d��H}f�A�a�[i=����TAj#a����#�NE�p0��_3G��\�U��U�h���Jw�4aH�R����'��5�^�&�ӄ�KG��*A;Kv��Ł�{�����j�$5��^�x�b&p
��ʕtu<e�,Fe݃Ƽ����w��KNN	�ފ�4�2�b���؏�hS*�DK�<�Q�L��)�<-r^X�_s��x����of2^���$@���^�a���ϵ��V��`���O�qÜ�}�5͉��Q�uhiY.�%\%�c�n&�`��[`�r��-��1�5V�[�N��
xz��!����������F·�G%_)���@j��*=���F��tg�۠��K����L_�?�� ڲ��]�z�c+@n_�v�ʭ7,_n���
:Ht�!��3$��L�*�%$[@VFu��+I�%���D�9b��vg8�!�Fa�A!?�s:Ѕ�J�*��"c%��Ҡ$���xwA� �kY�F�Ջ]�YE�?�`q��A)_s����U��)ݗ��Skh�B��M�P��f���(�N^4�]j�B>`f�r�>��F�f匌������=�ȑͶ�4K���w�K�H��t
���8W)2�Y֡��du�ѻ����I�*1$���c�����4�|q������;#� �3\�	����|���ξ���=��_�E�>��ō�z�����:s��
�� �1�VS$#����D���@���y:���i;�u4l��J/���)IS�Xr��C��Q��=�zG���|�]�g&�Q��A�%�����=�ߚ����X#'l5/�}6����.y:m�)���U�,��t�B���cŚ�$Հ긕�'�N��^�e/}����TzJm7l���B��D�����ܡ@����B�Ri�B�Br<�˛f��z)���'�GN�);,�0蠓b��R��Q��Z���N�m�t�?���c�?�,i2��!q�#.��`P���5�K�fc�«�0��ؤȈ�Ɵ
��W]@�[��E.ć�3��~*�]���W޳�O&/�-%!^��K����ؾ��#�+`�[��؉N֧J�?.M�%�J�Nz�� 4�p�����(o��J��7�p�~��<����&��?�Zxc�#��K���7j[	��B�Yj�7i��~ꢈ!
�/L& ���Jw�ڭ�$��̟���"����'n���sp�(�pӂ���lkH:.]��s;?�<���"��o���B"`\�+�;6���"�������z���H��o][�A�y�~��'�>�>~�	R�ae|NK�0]����
z�4��(�O��>#���E�#�~�4q�ښK�_��mDƜ�{t�sCZm��u��.h��C]��q�^j��D(\+�8?+�,P�t +�2��So�oFa
�~���	���>�%	�`��Z�M3�#1]t�b�����5�q6�E�埭�����#�؇�a-锽���xG-��}���k5R��s�XG�eZ�Nu�s�;i��Yȸup��:B%%�����i��WX+'��4m.�f?�o�t�ĩĄ���������n������q;�ap�O�+�OyN{��2���-tN���цk�i��I	��}�U�Ϳ�WE�)�?� �e���MT��A�c_9�]�8�:oV t%@��u��EPH��j�3�D�9���a؄��?������8�e�*���SRJ|�/�Cbx6j��,���Zj��I߂5s#)&�XrB4��\�H�S�k��}��>����&�v@���=����d9ᗏ�Y���t��#���ʢ+6�>��~U�Rٓ��JN>�AUB{��R�=�$e�K�Os���1��#m��xG��P����: �������P�SL(�a��S[`F��Q�0ƞG��#��`Hۉl�K�o4ہ��m�h{��������ə�k�d�@���9����k�!�ԫF�|���fK��1�u��j�tV����}�rn+��'Ud��1����J$or�[��{7�ʾ�L��Ȅ�+
:̹�bj0/�J�,4:ַ�z�6��/LTc�f݀�!J�7����9�1�"�Pn>��PD���[$�`�o���ȱS64�vr��9xp	*�}""vy�g���ܩ�}	�����������k���S�9U�F�r��8|%}e���)�WE8W�����A����\�fO�:���* ݢWX�o.�$&�w�}�D"��A2�?�1g�#�3.r����H���w6Bހhx �=^��&�z���JP��M6i�����++p��vB�&�o�gD�$�Ʃ�7��k͔��7�l1\+�=�/b�>�Y�+0�TS���]�H�� Yk��4凌�dӿ5��7LOPc�R��@8볟��UO*MD����k�7�3�	;�'��W������Ⴞ�����"�3g��hWL���9p�v�W ������q���C)��Q��9n@�������/!�Ȱ,T��ֆ��)���]Qb25j��� �*���`���S��W�Vح:�֙��Ke��L��"�iO�Sz����^�'E`@1�r����t_���w[����u^���T�P}���)Ơ�Jl榛&n5]M;!�b�X��tYE4+-�]���a�_�Ax�ew��5�c	:
�Ąƞ��|��B��	�V]��p�ن��/V����W8����)���Q*U?�k��M|���A���� Gt��^�d��Aa���Ĺ�@�@�|�ӫ�Ǘ��b^��~Ԙ�j���r�Лw�ǘ,�4���)�b��^���~�w�{�T:Q��E� �GA��΀�"2j���C��R20z�!(a_�3���Zb!Dࣔ��D᎘�?>D�>�v�`��I�&�B}���+�����X
���v�2
St\�9p{���V�o|��-'�.���� _�cF�3J��l�gY��òI�D��֤N���wDnw�3_l��G��$+���wZ���ϟ���&����?󤄰\"�1hU8�Lk姈���=�3x
�|nC�im�j"��&j�,_�,3�+m����&���	%��{zǼ�	X���EH�I������ %.48dG����&�X�wX���GH�Ӡ�P���}��$ܞC���7)��2�a6٧{����ۖ�_|� 6
j���\�^�iyO�=�����O���hWĉ=��f���D��,�?�HJ�В��U�Vd�W�o�}S��.]E�%~ ՀŚ(TY�c�I��}��3yPc� �$�63of�cNR�ߠ�­R�I|�E��ٝX"Ƥl�Ŀ옎h.|
ƒ���ATڴ~}v��Ƚ�J�h�)��ְa������e.p�2}\���U�r���P��=�7DMbL��1�ML,jbtX�V�@��#\����@#�=R*�9c�J�r~�)�i�'���vb��i~e��eW��@&�C"�c?��D:4l��y5��+�����s�L%g�T�Ob����H�_��%��B���g���_��GW��>pD��ˎ�h�gok{�������
w��~g�����t#�U07��ӿˮ3���y�e,Fq��"��Ǡ�a�o��k�<�?=>���]*����>"|�{���ź���Q�T^j�Y�6"�@��k4OѨ�GL�����U�f.���*�$X��+?���d\p��Qka_����(թ�o��Sr<�Z_���8��FN��'�rB�D�4[��g��2j/�6���etiQ�����r�l*��4�3/�����Ab�y��ѮAo]���_�\�v�XC?MF	�J�6Aɿ�4ž��$�Hճ��6[���!�S���p��l�Q��R���g���IW��}?r��-&SF]�������*���<c�y��@�p�l��û�z�4L5C�_����� +Y٧��#�Cn��	���7~vM�x<��]F��aw�4�>-�Hϲ��c�� �B�@|Tn�*�O�������-j��I���謁���'��	���u{�X��7���� ���!m�Z��	f��2��d	a��bݼj��8֐7���+���k��LY�g���Y+!��z��?C�>ӛ\�+�{F��܅����nB�_����=����&�bsC��ǤZS_�%���Eס�lk*������yF�`�Rw�<֡��R&�;�z���U5J�x��a��a�����MG���]yC̖����n7�<Z9����WFs�`L#���`╳�	{xQ��	3�Їnȕ�QI9�PUM��p���il�/�Ft��^��i+�=���U�z;ޢ���]s��0���3�P���Մ}zM�F9�{ӭ^������P.)��Z�[ޜw��|d����g͐c�萢�	<zR���Z�X4���bp���U��݃Ѱ��^��r��H8�zB��5	#u9�T�*}�	�ܱ&�O<�i��s-y�t��S#3���mBil_=i��~}qu�ھ$�'4��z�����lcy���ی��-���SMy� 1*�Tw��\��_��fp
�� �N���P�$��*�̫�5��/�^<��8�3v���֢�da�j�j��}P>��~w���"��.z�HCY �����1У�}�^�L2�l����\���΀�#g�9j�����!�|G~��B��Ł�0)�V���@�ojB��7�ڝ_of�����坶��%���8u�w��a3Y�k�~/f-c�k��o��
;AP�r���sԭ���+�n�͹��*�!��t�ѥ��Te�P�޸ǐJo�y3s2Q G=��;�Y��i�[{:K�11�ǩ�,�Q�]�w,u*Q!���̗u�4�]]+��x��Vvay�I�҃�b]��;^�C�G}�����Z�
�p�/[X��ME�<B�[���:,<����φ�V�Ϙ+pc�߮�ڔ������Dv��O��d��1�M�;�T�x��A���2�8A�����,��r��%�+Q�H�]u���Cko�|z�����j�H~ɢz�q*3&��H8cc&�jH	���[��dF�e?��}/�>��Bx���=�Ϸ�A�/���^K��k�i�>{��B;�%)�.��~����KM���8��VF؛^�K	��}�*��pvHL�5�S���>g�`�.�9�r���"�8�n�R��H5UO���<
ڗA�Mr�vW}�_��1��B��/d%���[��qZ/��-M���6L��ori��|�4�	y��˕T��!ֲU�$�=�	���r.V��D%T����u7��qE��-�����b�ܜ����)�V�m��s�4?9H�*�����o"(�{�W�����h鱩7&��ɵ���2�2P�����t��i<��P�}{5BQ)u�('̫�������9�b�e%;(����9�n]b��(�r�܏��¤0 ��7��g�t3���1���邒uP��BR��^Q�|�|��c�E�=Z擶��Y�B��##��$��L�̀�@c]אv�T�C|�KOJBnV���G��o��W@)K1��������.��4�HUh/���E�ή�1����H�J���ʘ�>��(�q!�����=�k1ު��O�	��<���jx�.��>!����a�i��Uh����F����PU��h����_����֙�90RC�~�L���۲��L���S�XW1Z�kh�FZtyB�Ȩ�:bX�{ve���E>{ؔ����̗m�U���S�o�=ǐ��,�߱P�Y�����O�HR^�+AT�]�9\>U8!�t�N�Vt��eG�<I�A����.���^#�O��^r��z�GQ֧����6��Ϛ#� ��Xu6-$���=љ�7(�^��SP���j}�������+��!�@3dpG��$&�,���ݯܴm�P걍=�����:C��m~U8[�M����~�A��f��1Y�C�*j/���QK�}�[�ϩ���ɸ,��9�$c�h-V����DX�I�@y QZ)�ϟa��� \z~2)�9f(
&�i�������x�h��I��Ü㦴n�}I�@��J�d��S�^���w�З�;��2�~��x(��1v
�Y~��|,o�l,!a���Ȣs�c����J#<}�����B���������N�����? �zk�%M��D2?v��V�⺜�1*�5R?�C.�'}D("9R��U����H!�s���+�����R�P���(3I�Y�5lU\� �'����㐆Ѯ]�!/_Z�n�������U
!�3�Y � �Nev}��,�r����2j`Q��c��,�䐽�'կ��ΐ�%� �Zz,��V�AK���\,*D��6��j��,k�^FΜ��&��^�#�Y��.�SdpMP����`p�$�q=˭���i�����~�=f�!FREo�*�nn�*mm|�i�s�z��)����C%��$n��$���H0*�<��e�B��VCU�[b�+��x���BA��h�� ��^�尓�S��ȊRq#�De�T��m4��^��߼��2)�6�!��ԏK�� \@pQa�ޕ��Ip��(��YA�Fs�q<\��8�s�B+�j������'yEW�j׃?��5�̣��c��e( ��c���/yG����t��Bb�#]h��;�H�����:��(Y��pW
X��t�c��Z����MkN��!8���5^ep6�}_�����Zq�T�o#��jB�b-�!��-�:����F�X�A9Pz16���+�f�M�"�1\TAwx̲����fg���f��b�ï��8�$�8����~��g'�]2��R��>�%�������gL�'� $�z�v�����P�@}z��>s|ܝb��)�U��PP���G�y`F��ۺ��vh;��V�q�֞$�N�[�Snr70��`��xfy�[��5�|�?���"%��F �;��� �U���Tb�����c��4k���bҴ��7��a�e  �9��;�*�6�|������l๱b�ܦ��z��O?�b0F�?,��NA�u(�C`�)/��O�>}ѤP��*z��D|	�9�r2�- �2u����V"��&uؼ�v�R��lMBL�'�A�_��q༫[�f���r�٥V:U�Z9_i#:z�kB�H�0��Nbտ�/�pt�f��ި�X(Ni�i�m`�T�A��6=���)��#�?���y��[�A��P'����+�O�>���h6ɖȏ��z��],�f΍�M�ELܨdj �[� M�PZ�e��
Sͩ~����K�������ֺ�H���/�`������@V0]�z*��nV���?p�������=�vֆ�z�-�&�/o{��:f��X��'�J{fץ�ꦧ���� :ɏ�^	�&M�_�S�5�Ж4D�Ҝ���N��5��SL<V�j��-���6ĸ,��zw�i}��O@	�/]߼�=ٽ�}����ez�y��@�ǫ���)�r��m1�	S���������3Y��z:o`�ȸTӦDs�U@��0�C����N�|�ը&Pl��>٣����ﱡ�U�@���XK�^~.���ڽ��̰P�^��`]mO�LY_ON?�d�=�x�^ڰ��j�ţ7n�_�jK�j����#����C���(�W�V:8`������xr���5��?)���e+��lI�|s�W��č��WᏰG�(P��5k�g����GJ�!��҄�?@��%Py��[.��������i.s)�O�s�${������\�K�s��"Ѹ��. ϭl�>l/	
��|����U?��ʮY��57�sүY����\�9�Q�^��ݠB���ַ����H�:���dˊ�� X���5m��e��+4ݪ�+��U��:��QW�Zq�	Y8tb҆ FZ�~W�pR%���%y�()�X�1uyri
;�u�*|����'WH��i�I��9z���q�"Z�Ԫ�Ê�@Ҏ�E���l�(r~�����M#a����E�.�m�p�����+�K�L�u|'c�;�
t&!Z�gO.I�C�d��H������7�M��(����$�]J���*�l�~Pڞ�zC�(���s��Bkx�KOK�ל�x�=�A��3�Pԛ\WS����u�����|Ի����
�� ���oFm2<I���؀z�����T�m7�σb�}5T����O��졥yw���d�|�C�1o!oy��kj�q1���U'jٟ9�X�V�^��fF��6m�4g�>0�H�g�m֋�/Y�&5E���[�^�2�﬋Ў�^Y�K#��ځ����İq�4��X�F����V�ZvY���ޞ9m��c�S��r�Kp��z;⭛���2���	M��+�iy�qb��DVLjT�]>���B���%�gR^g��N����B^�s�~dG��;!\��D��[�J�V^SK/E�z9�r��+O$�`+�AH/�:*�����E�1�-:J2f��[�Tu��&�N�$��� ����梹M��`I���[N_��i[C�ŉ𐺿�Yvw&$�̶_�RF߀�h���s��v�>� ��ґ�._��'��:7 ����]��W���2s�v�.&QX���T
)��,�<0�������p��E���1���?��S|3����H��V
^M*�pHqW��9���*�����F����Ă����yH4�Z�#��Zb�� �������U����lgi̡�-fu��@��&�mY�+�ů�!h��.��٧Us�R;*��f8?���,�]�}K�F��pᆐ�~7+�z�̙��'��IV�5I�t[�o<iD'������fg#tD�GR%�K��6�]��&@+�7=�X�x��٫R�k���e��
ں{Q��f��#��t��0�.��:�ِ��8����?D���#�����u0�D�fj���T�d��fˌU�O�ɺo�V�@�������sb�7�zJj��Æˁ��&k�x0����U|�Q�>�ߗk�V!��+~W�:)\#J���I�ޡ{^01��c�9)����E5T�t�s�ܑ����z�A�W�q������R�����=�� @���C��+�Ī�&KS9�e�>��5���@A_�rF�&�ȷ��[�^mʶ�16�B���..�t�ƺ����`Y;z쩼��̌yҍ�X@l��U�?X8�o�dX ��R5"z#ڔ��Zp�!����7B̓�����S��^pzvE�)�P-,}���L�7h�x9��".��G�!���K� Ɏ͠U" ��	��4P�I �i6�d�x0��ڌ.�*j��>��-��;5m{H��ؐ<�����Z�w�T�E���Qnl�A�=�H�7W�^5D�0ҤK�����J,
Q�a����|�����^�.��T.K;�3���y%�M���s�o�*�Č+����3�
kK�6��o��"��1\l+��DDY��tX�J2�k�I=7��y����&y�~���GG�sB�E�}�����:���A�,�kZ��eV�1m�y]#����� ��DV��i���s� L�幼q�:86�,f�.��<�l�£�Y�V�Z��-4%�\��1X2�|��/�R���]�Ai�����
S$�q��y�Q����d�큛�g�ci"�&kid�E���485��T|i��Dj�K;�u��rKo癩5@��(�%/�{wV�܏���rH�f� �w:m �����1?o��cැ3��o�x��5�	�{�u�a)"���>Ln�`Z���c$��]�eui�f����;���E1:�$�^�s:���瀲��Fr�{t��i֍��\�V�#�K��ߞ=9?/�Sg�=�d����F���!���D"�Ǆ��7�U��Mȧ�B߷�E�l�;'³�M4�[N�넰�j��>�!/3=���l��qSlمPy��.��e��G�JG�Bo���
�qO����R��t��7�E
���Ŵ�_�X[�ղ�lt��q.��o�/��d��J��w#O��wa����$^�p��O���UH��m�^Ô/��đ����!S��S����Q������e��!f��Ƥ�m)�rA-u;�����r����)	�+�^���#�]��>Pa��z�Y	�����eJ����A�<�]�Px�Q��[�m�m���mdO� 5������H*���L]�A�{�p���?� �J'��>�8��.Yu(���iq�t<U.��"�3�. 'f6��Xr���T��E�z�Ɖ��)��ps�p�Νڡ_a�!���Po�\Z��Z�k�+Q�g��2
Ҷ�]nd��՛*7w���<�+ ��$Q��E�{�"#Y�C܁2������f A<[yI�B?F_����+�������ɤݞ�`D$��*�쫨��V�����(��nCD���U֌2�xx�����/Ti��4;r�_o�!�c`�8ax�,_��X"쩁��g���mѰ����I9Q~�-����;mե���|�~4S �u9`��n�J"K��������z�b��M��Vmb�3��X�����kM���Y�a&�H���Hɒ6�>�G�&�Kb-Y#���<�#ӓ�`oV=�E�u���|V_Dj�����9XV*?���k�	��ʌ�#�wVU�)mŸ�e�T"���z�`�	�|S�N����ֻ��8uN��{�,�w��s,�yH�\��"#��#g,��u�<U<? ���  ��sP�$�yI����"ƃ��=�\�R�c-�>���`_�fM�P~�F��Ym��?y�" 4���V��6ip�;<��ꛙu�[��%Iޯ{S�P�0t@��C��4^.�Ǎ�+�t�)M|�����y�7vOW��H�h��͑�o7��=_ĹP��0�#��8�����;z7��e����	��~7ɗ�u��r���D�ޙ�!7��qG��;��-G���d�A�q�^vm�!Ӄ��i�)���G����CgAz�m)�xm�B�D�O�o����pD=z��~I� ��	��Q�#ͨg�s�z�ϭS{��_�0�b@�mZ�?0k\M������D� I2�v\~#B���B� #�',S�2	�J7#�M�D�)FF
}6�2�v4�� ,�y�E�~��C�)�d/tDN��jt�
;p�Unr)���YfM�z�IT�M���%��f��N��Lչ|�b�@�fK�!Y`E�D�J����������W�J���/�=Y�po�gW6�Eèu.��%���6v��������s$׊s��5׿�i����1[1c�`���������.������Ӷއ5��\��^ߪ�@U�N#W���4΋�����n%�u���^�qu�X.���J�]i}�@@E�љ��嶏�8�r�1�_�t�JT���sw`]J�$��F*�J��%�� �%��1��H����%Z�]J}��o�Qx4�������o���6�O��#C���j���aG�L��ߧ���sa�C-���S�4�f�B���]#:R�|	1���쉈C�/l�)���ۯ�L�W���Γ���R�@A������>/��v�	���r.�ј4����N�2�$��_]��V�yD��=���d��}�������W6 ���;+qyfN>̤��'!�DN×o��]���Z�7�;ed���6P�͑�y.q+��B�ps*8��߶ft�RZ���3�C'����O���t�\a��y��U�
î_F�v���ZB��a�; ��|��������A��"�\���9�"��poG�T�:Q9��F[G�E2��<��0��j��T����P��pU��\��_�L^���jI����r����K�$�Q���*<���!x�VE��P�q˴�ȸL�y����ɭW9I:��2�����V�33nwj�Qz����ȹŷ.�z����s�D�~/�=��w�Y�9�8�-��yʘ�n_�0,������>ĵQ��c��fſ�-%i�<j�iq��3��ӣ�Z�!Z��6[479��]6Q�{{A��ߠ���o�8��d����{��}2cZ� *������5N��	ם���V�j3�s�������q9����b�E+�YY-�d��X����G�~|�2'oc��B��O|e���
�\�Ɗ�7	N����٦���֌���1&�*�c�uX���X!�KT��;_m��ɧ�*
��P�"qƄʽ��V�`V��S�G �&-�Z��O��-���~�^,�[%՘=���n#��(�3��Miޔ��MkT��
���g>FO�Ǥ�>���P�� ݔ�g����t�F���D��	x��ϓ�-����0F�E%Q����DTtU��H� ����%M��"!_����h`� Q���B�;;�&d=%mE����H��ˏ� ����ͳ�����',�Y���u6}��|�N�+=b^y�p
��JT��kC`<n��3�hi	f�I����lK��P�8�?k�S)$�oIb�:�t%U�T�t�*�ʆ)�KFdךC���9�_���,{�y�©�V쁚}ꊵ ��nf�jd'��[w���� RW)�{ʧ�C�;سb��y
*0�;��ě�{�x�5��N͙-\k{��9λ��4j�L@h��zY�����G/��h�b*�FpH�*�|��T`�PXs�-�6`|tH�H�e����ei�4��o�#@�u��򕆑)gvz�]n#i��B`��I���d�mr�u�Έ�ԭ�ֈ��1��:M�=��J�=�Ѕ�t;Y�|+����!����A53�W*��t 2-��,ϲ���L~�NL��[��cȶ�g�vd����By\"�=ʞ_�r���Z*��.��0����Ð�ُ��WF�@�?��'T��.h�h��>C� ����:{�a6��o4��4������ݻ�\��e��b��Ue#4�8	T�?���-����Oy�<,�;�F��6v��LSu.q���� ��Z����:wCW7�7߽8ǕLk,���t��}�{��2e�/�:kp�1�h9�=�Փ�K�c���{���c� �8�~��B����X޵D?�Bl�I�Z��6·_B��L0Eĝ~�X��"�4b+A"b��TbF���z͜wE��S-v���n�D�3���N��6x��sd�N����e�	Q��OD�م�I+�,Qt.�>E�����H�!�DT����="����Ѯ,@�Sb0��ֹ�#��\P����u�7�-���T���Q�ʴ�;����[Rx����S���E��P�Pi�x������l�O�֍.��v���w���������P-���A�;��"�:V��� IZ�������[��F�惾���ʓ�5O�FW	�X	�������?{P?����yN+
��%D2?RU�=,�~��Z�g�|�/�Ϛ�ݎ<Q������_�� ������_�%�V�V�����2�H�ʳ���wo���%��.�������$EY2�k��A"�
�cDD�ZG@�������߫��
��6�7��c@�y��q��Y ����В�[��G�-�z�e�.+5���,�K̗X��QHUu�!�A֐ް!>��r��D\�:�U�8�9|!x(G�]��>����b
�F5�@t��ٷD�Jj_f��l}�¾�/��n�EJ�1�A:aZ�-�:�Z��r G���{�y���I�Z�h~4�Ui՗a�#B���L�Fh�\W�H81/*&���8�]MA3A~_�D�S�[NFq�Va�@幊<{�"r�z?��bJ�Tm���^���`���bo�6R��±o]3hp/�sh�h?,b��g�M�A�68��h q�_E2��L��J
����-F�礻��v	*�,��'<J��|Z���p �l2x���i�k\���0�w�r��-!� �F�4?����5K��=W��D�Eo�s�h��ZM��V4����{e~g���T-�\�[7Z�w�_��>LW�z��ϻ�aQ��(st$����S+������֚�3ga +�6�ߊ@���E�-�wh&���YW��v��=L���p�����'��p��������z�Z���Xi�|0��B(&/t��]��hs[\�oH��kBOǂ�I63) �b�5��(�¦r�q�@���9��Bv�c|/���[��J��?P��	;�/�C�J��
�%K�A��YOod$��_��0��v���"�`۬r�]d�ޮ��%Y���Rw8Ӝɩ��G5��
�wT#+(�ggm��r)C�6��s�ܟQ�zl'D�s;Jr��ߩ�S+2@�-Y?^�d&���dwR+���B�_g%A��%�𵥬�������4�4���i��]��20Je�MrƟuNCV��3�B�8v�kY��V�� A�bօ�\��Z��|Pu�,«	bMϥ����7�e�$���=����߮G�&��H�����o�Dkj�:�̷^)�E�Sz�|�-��s'+�_$�O��4?����1����M��
��0ԓ؁c���ɯz���x ����iҭ���e՚ڶ��:#�E&��]���H���&�m6�31D"\�X3o�u~�g㵁�Z�@
�c��W.@h�'֕t^����4m��M��~���5��!{�ozN81G� <�za&s��M�͊1���Y�B2�A��򗿬�V8N.��>���C�10(Фߋ��fb�ɖ'�p�| ż�W�c7�u/�41����j��8��K~tm��hV�q��YRe <�d[���So���LH��.%���r���~��&�6���ץ��Bd~ĒȆ�$\#ɱ
��¼�����F?�7A2�������B�����5��YRN~�=��X���jQ���`2жғȆ�܄z������*迤Q:���H�����8�~����vg����!��;�Y�`z:��)��>��D��V�'cb)�U��8I��p����~{�aҬP�[������H �z��m��p"��<T$�]X� ��o�w�-���!�԰`�{�ɇ�9����윙U�9�:�͸���P�$�l�.��S�'�x�G'U�8xZ�^�.1�?J/�K�
yݷ���U�/�^E� �_��%�$T��V\,S�һ ,U���� ҟ.�3et��dm3����h�<�n����s��v��KboB>��p�L	L@��8�G�:wyVg�^�ʀ!�21F�,�Hb�G�x��J.��\����(1�]W�vI��j�$�`E+q��څ/��?/.���EHKR�<��߸��+�$��.�*���-@r8�Uj�ԇ@v�Q�z����R�ow����TCUҒ��,+k�.�-g�G�Y��	]�ˌ�}�t��������^�����W;�����Ȯ{�)�P�J(
o�u����?�@G29��Ժ��I��n���3jr��e�W#�Z��4JhW�D�(|I�N�I��G9����HZs��������	c��obbh�h�������6(�LS8��y����Q$����q9Z�ZR=��{��SE~�0?Ũ�t�3�[�-t�[=��x0�/���	������;\(���O-�9�]�XR>m�����KG`����RZ�*��ƨ��5���rc������[
�SN��&Շ�.�fo��K�sK{R�(|����K�X�4h\Q<*W��
}b��j����S���OV�V
�V����9bGt-�S�_!	1��,����Ɲ-����� �$��Bi)��,o�6m�%�S����� u@� �vFb��~h!�m�t��,��&"�'Z}�ܣ6��;5�����C�1���Z;W'�����'��FT��9} �H��	
脊���d_��	�X�T�����Y�xǶ��h��[�.�RD��ԍ|����ԧ��w��Elq-�j��K�Ir�~r�/*�z>_@�F�{��3��3d\$���=��iD�'ޮ_����K�~�L��g��X5�=�,����=�GH��/�3e�-��ټQ@�҆Uho���Y��\@otJg7�ˡ�fbp}�-t�\U�]�!����gx�|�l;��Dq��\�<�˥�~�*�A�Ċ[��z"���:�"�|���*�DH�^��#�d�!&X�`Bv ���?^�F�����r��9&&J����HZ,~�r:���1�9h\b�u�G��8�YY���6�zE˭�̭K���S� R�c'K��nI����d��:"=-H��^j���d7E��N�{� ���ay5-"W�~j{�.�q- �p_��������\�$̟�"JC�����w|�l�e���~��՘�J�����;�+@]9<	�̨�g�L�U��୴H���vl"������J^E�|3��_�#��3��F���5�1� �R%G��0���h+�`F\��?V� �a!����i����|�ͯL@� �դ�bb�RrY���2��»ʝ����M�Vi�bi��@Z�m� � �[7��{p|Fr&�e��RF�J7�=����A���mZG�� �/撹J��?�F�tlǘ���U8d)V�$W����/F&���X�I���E�;uϴZ'j#~��ޏe����(�pj�Q��;�&�#jMV�j���D�[����_e8�����6#y��7���2F���X��M:>��} ��CZm����Lª���`���� ?[D�ek>8�|����؛��>��S��7�g(�[���+a�V��`�[��:���Эz���Zt��^�K��U�P�StpYY�7��V�W<��f�#�W];�*N���,����Nڏ���(n1��C%��� �Z*R�w`>v?�:��	�H��}�a�JR>
����;Dd̗�a��L%F8� �(i\܎���dS����!���D��x����%djY��0�$�'��q���QJ����0���� �xt�:��I��Z�a�x�8%ř��EX�L�5{��W�C�{ƭ��y���,�6�o�M �5���H-9 H��'@|��W(Z���`^�ƆTX��w���;�(���/v��L�Z���G�d�$��c�C0G[���0y��N@����`	��/Ȋ�qHc��&y�����[w������E`��ю�v�S�:�*UMZo' �eM~�����By��"\����������u�%^� _�9��N��, ��8zW���#���}���iHA\�ƍ痎��?GT8�T����K	�A Ƭ�LE#횫#EK�=R�v4A��P­�Fn���^���i��E7cr�Q��;������|�;��'4ɍ:��3ac|�Ju�4�3��p4oi:��F>��cjSU�v;l�!<)�r��������6Z݁�^��#�*� QO��k�V�vl�R�b���	;����bw���}�8|#]R�z��ii�	`�S�)�n��U����x��Ǎ����1���D4�M���DA���W'�����L�EdN�7q�R4X/�����=y��k��c	�uAX
���&K�r=@jѱpqc�~���Y�Ԁ	Z�2υ�0�NGu��VF}�[n���@�[��㽆Ȧ��9��*�O�'�n�a��:}�Y��	V�)>.'-L�}4�K'2�G��ڳaH���?5�p-wSc���;��D���AD������Ϻ6����;�\RE����?���[��l���ح(,y�����i�g�ū)����鱝1����1y���|�[�G��%�����H(���0l·ͦ�[�����K|iH�p�9��P��!�������C
��I��r�4J��i�z��<l�F��#���Y%.���g��SWɣ���*@`y�iƆ~Z���=�V5p�����(��DO�ے���a���Tv��BQ�4�t4�.����v����Th�<yWr+��؟�����E�7؉���C�X0�=�J��ْ��4��c�P��k�l�VA���#lR��熲R.�d|J]���tO��I����=#�C���	ך���~w^��h����.K2*Y"�B�����qk<�m�3�����/�`��A��t���︳�X�V�M[dy�k$�W�q:?�7BM���`ǭ9M�߮��hj\���mu�>_��;������	�{/:��.�Rh$K��k#��!�lcgyh@�����V8%J٬ʥܷCo�2��v���
���?�5�'�����sLr�>`3�9�c�24��+K��7<L���,�"�Z�)L��8����,_uwC��#7�F�d,������\�vlIb|V�����V��*ُ�{�����H~�1�I�#�V�*&�����O޳��G���5���VM��n �pa�s�=\m{��g��.?]��Z�a�����8��6����q��W�F�MO*�T��ڶy���3n��d��u0�^
m�=~�����I��v}կ]9����<�`v��M��j�0�PL�v���m�WQP�{�ARc��(�b�>b��v��Jn��'�]�<�(�]y�u�ֻs��el2�8Ή��p�|�/��N�H4t�b�:F�k��[�~b,�>�]]�MAhS��)�QM������P�d�.Mg���Y�o@��*���C���{�v9��+]����F�Z>k��& ���h?bW�`�!��N��������Їf�t�1^;V	��)G��J"�bz5{�T �7�[4�ӵ��!���u�f��+û�a�͇oľFG3� ��D(g���f��DA�~�il�AHG�T�'�1q*�m��D���*�io�����4Ÿ�l�씎�	ed�a����-�l�f?�L�3�vz,]�	���[���NB�]�-U��U�L	���ی)}
޸$�����x�5��c��?ncY�	�5��3�������^E��1�Z�5�3ن*�)�Z�F�>،�bV+�Ҧ)�
�]mc��Ze{�. ���/����a�"L��;���ob��@�Q�d� �͐Js�����eޛݗt�O���ÄւX\�����t���}2�K�rA���?A� W�f�ޝ��q��ˮY����I�׏v��gˊ�!��7��q�N�X����`<ⲩ�?��Ak[У�ת�2�M�D�(Ɉ7��0[Ç1�-<μ��r�Q>4�>=�'вP��`B�zyJT���[u�Nb	�b�+KR��)�$%�"�W����Fkk�J�B��y��vu}��MȱNR_1U*�i����/�R��I�d�|��*]-��3�E�q���I#%7�c��#R��t��������0�+ j*�9�^������1��ڑk��@��T���
$e]f &A@����a��%�t.&�JZe�#�jYm�����,�穳]���.���f�S�4��I~�y�^}�ˀ:Bҗ�[6�F�	��AXN�ӳ�GP�>N���lR�\��`l�uZ3���F���E�x���w�ZB��T�ړ��f�9����N��v���+����g�=�|�/Aٗ+�.%|�X+��e5n����Ƒ���I$#�c]�W4��ܧ�vA5�h�f6��2�W������I�fz�Ac���:?��3l(>,6�ܮd`�R�ǣ�Z'���/�B�yn˔C�#�o�o��it��*�������WV4F�0���Y-�}e�������H!��ݩG�ֽ��u$�vƋ&��#ɯ����u� ڨ��P��La��[M��;�4ڲ�:�8�0cLv�����-2�(��B Z��x�?��N��S��ي��TCf���y���e0�mC_�3�ַ�Tx�"oњ�^`����������bJ@�mH��WB����e��r[*+O�E��0���A��1����m�`���5Q7i���}H���[��"��W��p9��G��zv[=D���Swn��S��B�뽮(�
rRf�������J,U�L�i��"�����;R�2k�s5s�؇�j���S���Y'\�Y�S߃d�e]���>�&Է*:��Պ������<R�v E�V�j���ʟ���*(�u�@����Ԛ9�G��q��ձY����y¢D�E��j;	�t:y���>��ŕ6�i�(`'펃{���=��X��a��c`g�{@�P������ۆ�4�f�A/������)���]�I�R��"e�Qn�D�<Ϋ���(���Jc��{z�����w�HU��󽗣p��̳��.6V�̍���W*��U�ĕk�Ze�Z@�c�>G�y�qpJ�y�ϭ>~F��N��EB�0V�L��v8�����[��3��y���gl�ǐ٧8vHbG����P#��C[jg��VsЪv�b��d�ܝr�g%�X|z,H<Jq5ߖ5`��~ۊk�L�$E�T�25�5$)�v��/�؆=b�&
!�[�\���m�ijm&>wI�13Q���2Vo.��`T���rLZ6��QX��j�U°K�s��8~+ɹ�������̄K����Eisf�ȑQ��)G�d-$3n��(sǂe�"`���B.��<�1 h �up��<;�XXѩn��"ilK���p�;s
��C��R�_/J�@zU3w�m qf7������(��Y��՘v�×+AK�0����9#f��p��oF`�q���� �E�6	:?��zw
4�a2v�u��ey������/*�1�X¬�*q��Zd��=G���&K��J������1h��R�>]*�%��N�($Q�j��u�s���HM��p�������c�v7$�Bo��<�}���A{:�8�r�Z�����g�����W�S<�Cu�g�O��Hi�޸�V��E�>KS���cU�Q¨��J9B<��i�b4�j�x�v��as��?J�!�&����_�;�br���ӻ�[�<���ߪ��wc`fB训H?�'�n �,u/"��	8��=>����۩A�^$��Ҹ*����ؿ �]�z=���z�ϿA��7���H�co�J'��M`=�F�  Rq�0V����@�R�K��)�4��|~ ���~kbډӢ���t%��?y���R��zQ�� ����9��u�>����;��X�u����t=���C�����G���D���FL
��!�4���W��j�rBr>����58��|����Ơz�NUg�3�;E���h;X2�r-���.���	�i��͟�0d��}���ޚ�TK1��K�m�Pv��x �3��f��z�) � mXy��#X#��Ѿ���D�%Z�~���v��~=f���@��.�n���FK
cu7k�e�q��T`����4��� ٛ �,�0�]H��.( #y����;���^sǬ��h#	ru�lvT|g$��y��i�؄#6�4��F�xCsW|߀	;<��B�jtu���)E�SXtv��XW��"�;=T�����U9U�OӼ��(,��õ}H�79�eM�FM�l�0>�Ǟ.��"��go�^vm,�!�g�p1��#BF�W��M���E�$�ۗf<�,2}���Chx`�8�j�3b� �QA��Qk�96�:-h]�
B��_�lu~�Ȋ��+5�TM��@N�ב�Զ�`�^��3�I��~�EL��ѪE���<�`����f��a,��l[{!d@���r�>�o��̕9_0���z�B�!-ϑ��A�*�������F�)��ˬ2��ϫ*!�I�����9���G�1*��v[�z>�\fӑ&��9�͒�O�/$ߛ�� �?�R����H>)Jw��t������.�"l%e�
$�r����~Ɨ)��k�P�Վx�I#3�_���. 8|�{�fG���p�Q�a���ik�#q���sV(3�uJ+c�9�	���T0%>���:�덣�ŀi:�<�|�>�� %[��Sc�X�N��7ݹ���v1%����	8�{{U��f�)u�`��!��1�F�sT@��+����s��f(��ubd��E��D�!�^ݟZ5�c��:OQ)'���u=���6���s���\��U(C�'8IR����=��L�O��{ϖ@�H�Be�E��o�X�:�u.�x��n�n�v�]�zA�R�E'�H�|���O	7?�@Z�8��q!l���ӯ��M�%��[�bQ '��Յ��*�9т�v��2hor��T'A�1�$�`Z{X�seH��oIFa�� x��.f�/յ܋��J,�7�A����x~�c�O����ѡ
sS�5	ۏ���dk�(�Ȥ�E���Nx	f��6�4�>H�_�J�����F��:�K�5;U|O����[�(]�j�%A;�{�`����r�<P$�\R���Rzvcg�/c�Q^��<�u�,)Ǹ⻁���Ov3�߁P3^�!��n^��k��%���0`��|!���;T���HÅi��y�����U#���&�<��[_[�L}w�,zg��|ᙡLP�E��Z�$o��A�ꕹ���1�_H�c�C|������1��E�.<���Z���R�����S�^E��6��6�`�0��F���uT�D�2�о>eVk��5W��~�0Ŗ�!��0���n��Q���Y�4f�,�W�)rܢ��Dp-,��(�u�R'�a�ꌷH�F��C�5_ةS	�ͅ���O����&�K@��"�>��=���f�
M�vZ��jD�+A~�9Ӝͽ���
����5��!^���2����}�lk�k����|��t���}?@^��yx���m����f;s{J��<���n�+�����?##���^j8,���`����iEYI��?'6X
1l��m��u���Q�r, %}��[}遌��e+$ДcȜ�ug϶��K+��k���z�7V>i����c3��@C.-�0���I}�}�Pw �z-C�-��ä`⻆qR�EɺW��݁��+F�`�ꩨP��0�H3Sՙ��[je��o�
u�5�ߒ;˔b��s��[��������P0^d9�v(2�>m(�l�$\�^%G����(ޏ�i%��fŎ��P
�=��8`߫��:WƉ��&�Kl`��lj��R�ү�SjS�����@Ubؙ;�-�p���d���▝Fh!)���{�fȏq��x�Fp���7�&!�ؽx�ԝ�$�	@�淽�Ɋ{.9��A�X���ŦƔǒ�R�[�K����9�8Z�MT�����[�E�.����%61��94@�'��PÎ=���b�b��EP�Xd�RΟ��<��}f����j;���=��L�0�ޒ%�L��}n�2R*�4^�bþ 5�`ߎ�5j6�H�r��z��2`�vB�{V�E��Ѽ"��'欣]�{�ڣ���׵�A�b0
Y�pd�Ġ��*�)��r`)�G���'�y�e�&.L	1,�9T���4�[�+^����2_~'�ΰ �F!�i�ֿH�L�./�UƇ_����w��BRr��^}���E�C�Ų�G�70�IqX+��+w�O�����v~�Td<Ȣ�����w�n�a�0|i��28�=�O880:��N1㮦C	��6�̣��cv_����bk'�0O
H@�ҏ>/��e�\������@̱�}v�kc�7�O<��o�*=����A&�����~�]�f4�x�{G�^n�/�k����F]�U���������m��9���P��u��� b�`�|ȼ�\���`�U�}j2���C����Q�:�j̏���1}� ��Q��������O>��!�էD�旔!�O��)�!O�ay��W�	��8�cq�Q#҂��EwFN�*q����H���&�RU��m�y��t$ �%�m�Y����#*(\,���q��I��v=A�(��ư��*����� �j�؉rC���D�vi.F!�h����*���H� W�
!l��bU�e h�"nW�Yw�e��a�A���0i�W��{2"���a^�tB�$��~���\x���$��u
:��>l+�BF��KZ|9���|�s�s���2�$��^Jϱ�ў��2��ځ;z�DSG�ӕI�����a���xO����:%��7t��%?kR�?���(�*ݣ(��4p��->y82T�i�$�F� yS*��?Ȇ3���cI%G_DT$�����|���Ȯ����M^�ެ��t��W��;f9ʿ 3'X�H.��d*�t/°��}�=�	�~�� ^H-�A��A@�l�+V��ڋ&����]��Tr`�Ye���*��pPF��x����oki==�A!���7�ǣ�;=�E���@���P�f���&[��/"�H�1M�j!F1*�@Z�_���:���!��:��R�
|��h��w�E�����ug��7r�> 됣Y��ة�?��t��Nb���a��7,��?UC[���	�g�3�,z ���|��z 3�M�_	L�]$�3���?�! 4���;GUj/��	�C�����-�]��aZ�-Y���^��,Kg0wv��;��g�,=�}�4����B�LZ�*���ޭ�۽��1� C��(��.#;�NǑ�Ā�}e����?R�v�>a�{1�*��o1��tM˓��#��#V+�C8�+B����`��g'' ��"�Q��N���`n������3#�����n���)3D�D��TXJ�R�>��<K����@Y<B�l�&E?�<WPC����
�2O�v�/K���9�`�
���~S Q��{]L���^ց�j,���:�~���90�����l���nW:��0}���S��4x�����7	c��b��J�'�f�LZ��_�jolW�@-�P��2f�@%��Vŵů�n�MV�e�A���(˅�$�u�?�Y/�p�§h�m��f�O>�f���*�ᾌ�s5i Ê���7Y$��[t��ӗ��n��˦�����?�����I�7%�9B�NΛ�*Rn~�G�:r���]z�я�e�XF�����]����yݦ�u3љ;6�;Hg����r����q]7Cܹ��B�U0�)�ke}4<>~)4L)�hҾ�pu��+��jއ��nI��E��X垳�Vߦ[?c�X�A5�S�<x�F��9�����tw�ߤ�3��9n�;�,��t֤��{�������{Fb0�%�# �/Qo��E(�`�::��3m`��Q�qⶤU�/�X/�� 2���� �+��$��a~��*Z�Ջ3�[�}��r8l?�5�VAX˗[��u��'�N��-t��Jt��Ê_����	����p���?�B(C�%b��-N�{3�x��َ9��_�q� <oI�{Wq���%50�*��>��b���p}�¯��Kwz����fRq��QCL@���c�U,ZcI��Z����B�pƢ}.F�}3�?�ߧA8_f>N�^�y� ?��K��KgB��Iu��@@���v�`r�l�$��� �pd��EI��wH����=8YMt����%��q '��$����Z�gU:��B�=�h�al�#~� P_�����/�t�+�ڔ�>����� ol�VQe��-_sE%�2'T�g�.������~��4|�DqE(����'d��:�_��ʮ�kb2�g?ۛ�|R���A��~Q6�����z&��F���d�j�6K�o�T�t1�= �#=�c���F��pqj�P��p��� i]����PB11�(L�1�oI69�e�f<���O���3g�f��Y�T
��=�j^���F����J��
�X��>ƙ��Ya�U؇���	����ņ��?�$�MA,+J�Y�q������qh%V�����|�?����[xwu^bB`�| L��*6u��] 5K'r]�J=���J纪�<}����-'���H���������s�||ԛ��
�(�z:�"�����E��fs�����1 ��W���c԰�	p��}1wl��t���9C�YKIm�0�1���u�-���57�����N��@5�F?���7�t1(q#ś?y��?�����ċ�E�'�:�Q�*�w��*A���!����R]�n)h|���am�U4� �&�Al]������l�_��ta�T�/7�(\]B���#q�9�A+�~�k�����P����ئ�+-�|s�H�������Z�{��
�<C��܎n�cW�$_�_�M��W�F��C�P����zƶ�;"��iI�J�Hz��c�(�޴���8nXVڍ-b(�W�y�^�h.Ĺ|��%���#�-�f��%L��{6n��K}�.W�{HO��
�s� �<\��f����vX�f�?�m;'��e䬬�2ZOT�J�Y�t�_�ZZ��"C��N7L[�	����C2�7B	d
MŲ�7:T��*�B���w�b�����1�;$�V�Ϙ��|+��p�u3͹'6n�X����{�@���r���G�0�8���g��g@gmꖟݜa%�郛�&��aK���cx  Azݬ,�[�T�=h�C���RH�B�N���F kb�rGi�(���w�E2���kn'�� �Цc*���e�S�f�?|�*��
��~��K;�kùc/Y�
q�x��QP2���Gj*�Qz�8Mz�%~�շ�>�ĠD�
����eŁE����eUu؈���L�7�����Pv��Md|6Ϋ���9éDe��i^r�����e
���8��i�'Jr�]`��_V�\UM9{i��z����#ć､�=���h��HQ��ޱ�րPeZ����K���q@}fl�7��m��=LAf9�1]���C�!d�I�����,$^���Y�����|���|�9gh�V��f�O���.��~���we�N��&���HQv�Kq���\&b[��9^{(S"�#��{�ׇk�[)=�Ԅ�Fgچ�/��omk����|� ��YOQ��α! ��
��=��\�ۚ���M��6��6�r�^���͈��)�tԪ��UW�9z�k�"n���&"�%{�\,h���I��u��kK��l`^��/�J�}[�rJN@{�N� Y>^��0&��:�vuD��3��V��{h.�i̞D�2(��'<)��1�;g$�O�+����g��S��w�#� ��k���?S�xʃ>��:E��p+������L�����p���}���2��x��O	[�Ϝ��r��F�W�ɞ�j�nP�������"���X�,??P�;�Í2'�ԥ�|���XK筓��>�֕h�&LLҙW����dH���g�UԄX%^��:f��)�9�F�EY�H��L���<�Z�7�����`����~�=�/pq�4}DTK�r�F�=;�I4)�Jk)Wew�{���4����LC*��l��w��u�v#���`�@KyFA�K�~��v���I���ݍ4��_��Y�cQuK�V��;Zv|���A��<vjtc�C�����Ыݩ�)H�
�k'W�y�c}��ZjGb#W�0���T�-K����*�y*����C75 ��Ҷ���ܛcUyC��=�+��s�K��^[�q�RK[J�)E}��1 t����E*`�n"��"Lw�EF}���'��У�*!@����,$s�W�l��+!xV�/\"��[��g�o�96l���di�O�.����xI<��%}�:�(���L9�>MC,�Ln{,د�Kl�ޣu �,�j:����� )��0�M�N�*N�5F:;DX���_V*B�O.�s�Ls<��J��t���ҟ7�d�����v~��	���y�=�\�s[N���Ӕ,�Z�[��(o*�^�+>J/`�l-�u89���>k��(��tv�u��
���Ƞ��wb�8"ݘ�'�)Ѳ�|B�M�P>M'P1�q�e��A*�+�0J��(�0�@05�:z9�Xe�����I\t���,�Y�
a1E�ǶmS�;.�?�63��s+��/���xX��AzY�Յ0_E�3`w�/��G�	fQ��HQ7��#6���Zͱ̭Z�w"b�����a�V~������ImԀ`>}���ư��l�ZdF�������US)W]�u��S^禙�����| ����#7k�:֔
�@'���i�q�;���M��-�;=nU����?(/��ȕ����Uo]����85��F4k{gCU1�~�W��/9���gv]�y�A��5����/�b,!R 2KЕ)��K!
r�����F_]�)������f�u�1ě��M?��U<�b�5�2�!�]in<8�|~-���(dk�;R�\�HT�[.v����^���%�ABN��!�������g���%6?�=_څ�g��6/O\��+��K�)� 1\�'��s��|��"��~%��p����O,7����a-f�ׄ:�*��v�-������,�&7�2 ��ܞ�s1m�\h>b�0�i�x���o�1��3�l�Aע��~���$��X�\�O\��!	`$q����T�!0UV�]�A�S!;B�*���m��^�<a=i��k��/��>�,W��{9��-!������,��˒���Z���j̾Ð5Ujf�k/o�[�^�>>��/����Z҃��>�;x�FV-A=_��kC̻m���kQ���/�uZK�ʤ��Y J�>ql��:
�-����D�j8ɖߛ�
."}����=�.��V��}���YE!����Z�+�uMv�֓�sdD�{���<v%h�)9W�$�WV��a�t��g���+5A[q2W����{�Ԩ��~��yo+��n��c�m��A|�Є�$b�]��m�$�/��$`��պrIg�-$:"<��{���΂)�f�[ǋ,˵Rtr�K���l��l�[�q�f�+9c��9[��jt�G�D�X׾�ѥ��y�9E[Ǐ%"zZU��ei8V�cUȮ"]�jtxcUf��� ��ա�S{��	���C����L
���DO�J�8�a|�;L}L�B"�c����-�\\.��z�o��w��SG>F$���s���}N� ���(�!���L��q�wwq�+΅3},�)�蜗�-&b�S�O���=L&&�-�;�'�/�,OH}%�b")�J@nc�8w�R`��w@|���\#@�P��rGj��S���r8�I@<f$�(����b�y�A3�ŏ�egP:��ɢI � �ŏ��]��h{�-�AX���4S�����Cn/2��V�&������c]V��Yce�8�,��BI�r��AQ��ft��'���/�.�"�W@{�S�>6-�w���}�B�>��!S],zO�V�����~�O�a���$#�J���W+�!�A��)ol�[H~lM��k������^�G�05~����t�S���<����
|��z�~�I�Q)�s�?�_=a˘ʽ[�_�֍�jΣ_��Rfv�ma��")��R�q}`V4W%���a�m���OM��L��\�qRn�*�������n$���5c���OR�[�w1
za	�d�KۺoE1���t�@4��A����TS4 �������5RYW� (��m��槲�^��j�&.6�!nĽ�|XQȹ�\���w����r����U��Z"��&�Bz�:S5�Ux\_�I���@��vF��L㩫1��r=��G�r��>tPq[W���ym�l� �|bI���J��a`ZD���Uk|Z#�O<�¢[���^=dO/���[�v���"{�p� �	f�=P�O�ц�q	VG��6Z}��#̂kX��(�-@�a+נnLR�]�k�h��Wg?���*��0���(�=��n�R3_�%lW3�� m�?57y�²f��LVӈ�}�]�<�cw�%f�]Mˆ^�ܖİ������v�x9��l���f�&�,!c��`?�lpr�Ľ�ebU�4]wp���!�̛I��������6C�u��j�h�a�-�Kr��^��'>��X��uhcum(=~�d�vm瀪�5�^<�o���W,�G�?�l�X�(�\[%_L�v�缒�>6�5yʻM��	�-��
�*>�n[P�cJٌ������KG�D�|��a�&,ӷ��>9�$�)	3..`�&ߪɬW��׹����V�WKUse2f-�^å;�t�ӳh0MH@��v��o��->Vp���D@p���ޙ/�w�#pHy�ђa��vNF����`�D�w�/;49�C	�t�E�ę��_���g?CvQC�sM$/p�O�:g�=
��gV�qD��^�ܢ4�����Z��g�۱ȠY�kc��<���ӧ_kU����$��^Gq-��s��X�{�N�����`��z�;��.xh����+)�LÁ�&1:׶�A| H�b�y@0��Lb0�K���������d���W�KˀD����ջ&���
��d�?a�5�|!��z�]4�JJ��(��p��`������Inx,���-���λ��X���d&�bS���vn��JoAi"�ܞ��(���w���V�Ft	�+6ڦ���:�2}�O!��!R⡰Lܪ�ʗd3�ԫ�Nɲ�%���$�.>)�bt3lކ����{�ц�j���v
��h�c�5^;�����-����~��B��jm�λo�Y6s����i�#�{�X2�^�Uy	s�H��}b��6��[uo�2g6c���6$D�q)�:S����y}�؅ϳ��{�<�.�\��ɪrG4~T�C�B2ف�K���3�ğ=�p�P9�	�	�� C��=������?��:��7B}R}v��J ��4ӣy�q��kz�8%�I���-����ADƧA���k�3�}�=����)�8k&�����E�arF#�P���‷�mǤ�Ł�a_�`fVqV�f������ �p��}͵A�з�U=� �|(Ҏ�M1*�=ƛd�v�P����4�AS�@v��\|KD\�iP����Λ'�؇_M0��2n�	ł{�z?��#��~~t�y���K_e��0��DU
���1J����`�r���W
��dVǇ�.�sL
�N����`�%����"Pf�{�L�1�h�n��f��
%W�j2�~��0�M�>|��ʦ ���E�+%R I��yX�2(�Ơ���\V
[�xk�RAaƆ��3X�8C#���!��y&ީ.;c��L_��O���3��3�5=v����v�S?��F�;K�sc-%(q���+N�n"D����`���mC'^fCcy��W�ӎ�(� ����8���:2�}��[\H�`W�{� ���^��F-��x0��tog�R����?����Pۧ�-ܵ��X?ͦ��4��<�f���F�Q�0C4A�c�*��kXȂ��r��BC,�E�66oN�U���Z&�8]�R5����������`�-�K��~E�a&��V�U.`9�����8.�}�U��p��`
-�Ga�q
&�;�?n[D��1��޺dXf���'l��\Y֮�~�$)�`u�� �o�l���� ���}ir_�,2���w���as�]�A��mϾp8s욟��k{^$�a�B�tiq�т��٨#��$���EFl(Yj�s��ɘ
�3�[�E�i�g��լ)��$i�Q�d���_?���7��g-g���چ0�}7��l@�Y�����ۡLk�(�q�\���,���x�
?h��E���F����18ʲA���=$���*�fLmf�k��6�%/�y�i�W�/�=���շ����}!�0A�5��o%G� m�|*N���<���o��x��#zY�wl�aq�Ҍ�P�]Z�M���A����\/��b3����4�5]M��kӐ
�{<���ª�s$�|����yx8��n�팊��k7�H��)���%L�.�x�O^qE���z��1�]�'�b<�������"�v���m��T>
�P��M\��V��7Ej�("hF�P��O��E�	uF\�d	����:FL�%��*���y��06MO�O�I��V�k�r�4�@	���9}u���N��9ѡ�"�;���e��}+,!�шEs�;��af�w�R��E����*߀�`��Y�u�`��{#��<�O\��{�������J4�I��֏
�a�膄5�ދ�� +n���n}��4�����Dpz�j9��G��LB�
�&�ؕ΃���x.>�><�z�;Dʨ��=q�X� (��֮�Ĳb�!Er�����=��'�Gˁͨ�CB kl�	Ba�tn�V����4ъn��9e'��D�J@��:��Մ���&�_��{��biHj�U�W��!GNke�)��D�[�T4�ܐ�F�D�\rS��OH}@�e�Z�;��.fbb�Җ�����wbK��d6c3M��y��7H�LӸ��j/�X�&�Af��y�Q ����c�Z1fpf�ﾤ��b�M(��3D����i5���A�7�P �U�ȑ�~���Dt���i�A�h�f�����cfk))��r����)#��$�K�����K奁P�
)����~�]��*�c�C�!��kN4���Iz�|��L��~�z 6��Ǝ��/w��15���'��9X?�S�ML��̯�T�9�OR�M#�7�f�U�l�u�����y�E�G�����5@j�6?�؟Y �Бv
8������%����2YFe6��Ht�$��\@�A�R�,�Ap?�L�#����_A���>0�4 ~�H��o�h�Z;�]���zN��疶��r����^�T���VUg �>}�A-�(��/�F�<��L���v����`��@ n ��t���I�k�3��t	cCv���R.�P1�6:���k�I��E�	�X��E)
qF�#����](N���������(�5h�ކ�PT���8�ջ~1��/24��q���9;<6歑�g3�^@[]}��ot� �P�R�)����_Ǆ=w��eL=x���B�3/L�a���B�"�����-	G)�[��ܱB�
���=N�((�.�U)�VQ�LD�g���Fv���=�[�};U�T7.�檉�M��z7R�l3>�C2�Ea"M(b�T�ϫ�.��'t��ՠ�\:J�;�+!�F����Q $��وS��H�8���a��=��? �Nv��ۑr�母FV�u�S5c0��S���K�����s���u)��n&�N;'r���)�!Mt�����U���1����[�mX�?�؇�[�_��Qo��U�<b>=��8�Z���	xW��!-�iD�G�>q��.)��З+����d�����ч)�sP�s��`i����[^ȘfW9��-U܃s�H������\��b�'c�)܊��=7>6|��֖�����hv��mE�����*.�7�o?�X�s3H{B��Y��^�Q�͟7eVFh�J[��²�_`�����������u]�p�v�05���+/����5 ñKu���39%n��]��?���U���C���4���Gs����:��fFU���ވ�`L�稴��MGF����I5D�|��S�����AfA5"�b�B*4R�u�8�22"��ڶ��aޒ��V>;tK���2��{�A�9���\Z aUdv3��zs��"Wh}=�HD-��"��~1wT��&�U�j�ggK�+�!� {*�Ȟ���$�}��8�ɉ2O��m��!�V�	���<֚]K��3���ؔb��&��Y�� ܞ�Fb�EnK��.ڕ���lx7��2M3�\L<�p���xy�JS~R-_i��}z�%�s{JM��<B3��g��,�*�x�T�#�{!^�Aq�J���*�*�����K�O�}�3��p���\���=�L��m�����S���7�+�3%�R��@%Qq��K.5��-�ڼcw���?��;�S�j-n]�����)�`��xπ���˳MRjƫ�+c6���sT��#�ԝ���%�Y�a\����6ՠ`��S&�1�߱��?׾tVs��� m���5nE-qu���B��WV������9�#Pp={d�6f"�Q�?�����}P���!����sZN�V�����C�����}t1Mj���.�j�N����h�����IjV2EB���MfnL�K��B��-Ѧ�L��u���g�*��!9��n��阈u�4w\W96�d�e+s�'�c��FF@�
��Zv�7V��O踚Ѷ�"��U�ϰ��x�KI�Rx��2��@���F-�N����� ���&�jl�,Ž<Z��`���Ӵ;`�cp`I��`�)<ܩ��f�k���*���ߞ��p,(�u5��=Uo�;�܏il�2�`i��Д3om��-<�����;�X��HU 4���'+��c��'��v�qK���L/|Z[��x"��9����J�nP9�(z7��&��(�]e��0�~\�;�1H��>��c]��7�ޫ7:I�S��de�*��xG(	�78"-�G��0\�<�ďI����K}�m�5I3ъ&���AKO���D��v4B��̀�c����bm]�]v�#<%��	�<TL�*M���ֶ3:�De1gB��}�R�N��";���/hhfY���� ��8��BbI��.�����7�vs�f㐼9j��m�.�Q�Q�5o��k^����^{���ˆ�( ^�:I��o�	��V� RQ103@�6��M��tݼ� ��� ��v��78��ʰm��~8�Sv���γ���7F�����6a��MI	�dNm[b���qo� >"s�(}b��I}�J�i�v���e|���QϏ8)M���d�f�R�[-�#���`h0�ό�%�����)�����Z*/���ڒ�O�b�~q:� y��_��OZ�>r��:��ϡ��z�j̨�d�s�GH*�>-A�R�ZVuEdq!a۶��-9�s�w�5z��|�p-�}���'�R" ��M���k��[,D-��k��?�1�P5��з�^�u��B�[�n�g��k��xn�;�H�X�7�?�z��B}��::������S��5��iq� ��G2���>��|���T��4���<�J�R$�;�gBa��qc��=��>)nD��º�� n�xǗM8��pSB#��	�I+��,G_������5�b����JG9zZh��ت��6¾����H����-��� �t�ް����#:��W}*An)E�o��c��Hq�*����N�^*Ю9.��ƠB�A�V��8z%��}Å��r���Aە�r���5�?��� ��7�0Q�A�(�JG��ںG(�I��.J���d	ƶn�.���}%Ҷ�{�d���X�jR��KOlv�B��OD��� aAFg ���u��ĥ�͢�*�";�,�:������\pB��WX���S��0���7>M��.]�>�)ýe��p��;�<PXȵQ�0!�|]�D
i��� ���f�P�̋�˹Q0�ݎp�r��� ��vV�(Q-�h.������n��}nٟc��Lw嶼��S~4��e'��H��ü�pl ��|F�kpK�|\��n�6o��{5uQ^�:�����O�#�گ.�{�5;R�" ���_�2�`�r�B��G�:�2y���Y�˰��x'��у�����q�kh-m{���Kr�jgӖ����/�(��9��:��F�s��V%=���O�`�5�H�S9��!�7�.S\f���Y�0' "���3sx�e	EeS��e0�cv���t�+��#�� �ڵ��4�>�K�L��٧�T���8��$�����E�*�/�93�p�쉕 ��oz�b]E����#D_���Q�\S��&Y$r|�e�
z؋p9Qgh��kO�=�N�H9�m���ÁG�ʿ��=�e�:�K�*��v�Y�b��
�/��y��dj�ɞ�hBH���agxX�͉? BJ!#���C�}��HRN���B�&T9��mG�>[�)���j��-0�E���@^Ej�SJ�Q�O��^)����yTӶX��`�\�k��� �S�V��I��5@��)k�+��-*�-��$�8�)q��N�D9;�w��\z�ռ�Ƅ�m�����/kb�
��H9�3��|��=��Z1��(�9�fV���g����q���7O/��k�Y}�m�b��ǮH܂%�:�.�<hX7��)}׵�e�mO��J��X9��������ϟ<�����@�ASa}�a�܊�?�a�u����%��w��ݺ�aO7^e ���Pk,�i��9�&+��:�q}n�\h�"�H�K�����R���G�6P쎺N����ߪ�آB��{'O0�@��K�M��_�0iR�:��g�?�+7�K�f��B��/�%&�m��̱藁��:��ـq<,�I�h��T�uj	7�5 �y�@���/)�p�����4�n��|�S��S�%_��k����R�]`5�RyW-�{���N��C]�ڜob��)k�Z���Lw�ֿYe�D-ZԒ�J�{��m\%�	����eЊ�:~��ӿh��NI�wC4�]W�y�����S���k˷��(|p͹�ޔ�lk���^B#j�y������y.��)��,HjԘp��\����-&��fD>GIo��it��L$�P4G�1��k*db^m˗��A��]�����;%V�Y@�7:y�vT&�G�����~Bo�q��Bﲒv�jg�w{�'�x -; cF���+z��yNȅ��z��ָ�Ė�X�")�O�7���u<�LOii
��y�ŐaI���'��@U��nZ�$QY��A\�xA�&����4���N�6C}��;FEB׃o2vj�>G�5���i�Ջ�}�F�e��O���1�R:N�Q���@L��G$xk����a�ρ7/=�_�K��9_�CN�}��I|��*�uKTd�.0��0(�m ���*���!�C%�!da���؂�_�я,�:2!u�/4�����9�f#��#�t�m�g*��][���� w����Y�<�G	JًX�}���~�/�|�G��ʎ�����z�K��]��eŸ�Tvj�"�A���ȗ7�L��ٗ]Hb�$�K��������0�Tm�9�������um���J�\�i��xr�l?=Kw�@��>����oG;U�%�wߘE.5nʑ�^��De�AF��e�uu1q���ٺ� ���-��^���Z�Z�./�-����6I�Q�.T��Sfӈ]��	�S���j3�1�i����#�Ӈ��-���іۏ$�{��J	��8# _���D��Ī5KP ��S)ν�ޗ�N����sg%��aM2�#>�M,���؈���,]E������8e�t��I�����+џ(����;@���}r`�HW����1���\��I(��Q��iYk~����V_����X���ߌ�¿D��J��-�-8�'�n�u�Y�|�Cۈ������L`XE�f;T�p&muh�c�O�
��o�P�^�����Af����]��$�s0�GB�oR̖bD���h�,�=��	h��,����ɞ
�ƽU�I�pIC��"�!��uE�3�8�Ò���
)���#���׾�T���q:`=w���(aRT�H"6�.k,gr��q0�e��W�}Uw&�u7�7 0_��v^��;}1�@�"cNt�v5i(e&'s�O�k���>�$j�=[E�����n�\p��Nw��ZC;�^N�-ܽr�qXi�MحM\�"t~E>������3i��Iܫ��7 t_��a���͠���<h�!��TS:�J; µzi����	n?hR���eW���%ä{��&�/貍~��)B��4�6[����/zSb:��_�ճ�.96��D�R�]X��/Hi��(:,�]X�P�e;�kpz���F�'�A��&)�oåYE��-��f�s�x�u�$B����g�s�PS�� l:�.�.��ǅ��,-�2/�>d�*j�X�M�M�O�iO�Y1mG�B�%ο7��
v��� ��u}������S�,�\�Ra�����U�N1�Yƨ(V�9_�X���%���,r�,�7�q?�}Dҫ�ĵ��+N�8������~6G�+�����W��1t�5��.h�ܳ��&�m�e�l�u�:�q��o���G��#���[H����F��Ƣ̙:��&=<��-W����5J_�"#�0N �$��Kߴi�gt��r� "Ŀ;WH�B5��4��2��c7G��9T�k���[�4�7��vF��T�]��\�V�:s5BQ�OhD�!C�E�H�������}��J`$��8z�{ם�3�UW�ȆS�@��N'�=r�2���A��>k;Ե��v�*�����:R�����*,��eG?���%�����{��/ӳ�$ ^sW1�5���*��y�(�X��ߛ��8�3�A.ֻ��P��7��S���.�1�2#�f��_xj�Z?%L)K�z�o�57�eT�z���L�SW��O|ڌj K�h�yt�� -@�`��m3B���+����n^4���'�?���E����Z�?�ߠ�~��OU[j쁕r� 4�7JU,`��ɶ�{���Y/AQ�+��0��	W��!(xsf3�ʫ�Yp�S@��e��yg,�Ii�|��e8o�]�I$3����DI�X/���[�2�Q&O;A:�é�3@z���	t�աT�"�j�z2+��?���'�����q��>�	N�,aȀa�� �yB�̊׍��@��yS��S R��wT��imF�)�K�JIz��y�*�����=�`Áf4���h�d$����5�u��9�% U&*�-i&�͎bS�uF���|+K���B�6B>檛�N�nU���l��D���q�8�m�!Pä����.�e�j@���,�+]���?�5��`;՗
5
@�`l�;��Q�$��$r�@G9��s�D�>�LP@6���C!U�������ѓ{4��~�nW
��أ@:��N�W���w ��'�,hoU�<�3�q�ʐ�ZU����8�+=l//S{ȅm��ͤ��E��N������Q6�����\U�����������ŰD�2�;��"�k����z��5�����xS�,_����Y����T^����Nޔ�/�[�j�" �)ڱSR�1��:f+SƂ1cv��V3�b5g�2��jqY�YjJK�z;B������x��#,ҤWu����#��c	i���6���]� � u�c\-*���Ep�[C2.T%y��b�$z�?!��y�r$<G�4E#Ǜs�~�,��T
H�O! ���#Y�C���b����J��$W_qUO�zܶow��q�\����F�r�ˎ0�#i��D�I��{�Z�R��������J2��H��;U����r�nvi��&��~�̎��l���Sb_����pTS��°�#&[o��S��՛��_�3��i6�
����rf���Pqدˆ(�_�>NPP�����e��{_��4� ՚_do��V}] �Е^B�m̪A^$�.AQ�������t�I E:b�ɳ��Ȗ�����&������%9B�6�H�"�y���[�ͺ��;��5�9)�4��2� �����J��Ǫ@c�`u3Tr)�
��B�,ˀ��	�>L�͙����I��ܼ!a7=�m����b�;_7��P�K�ʦG�T�.?z�ڷɏ�0
����X��9��|os<N�)�{����H�5�w5GDԂ��W���I�A�.W�#���p
�oY���M���]�
�j�L��L#>,K̑C��I�8���P�l���;�V�LW4r��$��>��~{e^U���e�J�/�`�h��1qL�t�(��4P��YP(���&ՒP�)�1+�u;�1�̇[S^�=�B%l�Ԑ��eb����c/�V^8
zMg	nY������?�\`�Ѫ�ȏO3�"L�-���p[�۲����6،�U!�LbA��?�j���T��t���d��Sfe�#q�eq�>׮�TŬ)�q�$܍�/%*���B��Ii���>��R���29����ST󦊥D}(��ܶ��e���W�*L_W��G͟�W�����j�뗒Y��-P:u�u�o�ml�MMA��A�4i>������d^F�t�T�3���8�=��t}���B"��ٵ,ּl�Ax��bT��-���"��R̩�+ݜA���k(�"(�3B�\�ڵ�â	a�G�ݹvA,��-1�2���8�a�.�� � 1�
<դd��-������Y��$�D,���|kR^����,�_'+�x�{�����h�0�x����_#T��@�.��{��+1X�;ݮh�ȏ�Ӝ�n/�q�i��*KֹST�3*�6 %*�҈�����I��[m�7����٢�ǭ�H.���W�nvҁø���TK�2��
�L0����u�01\}�l���2���_E�p�!���&A�qj��^ƒ�w"�v▦�jp�x>�gͷ����<��׹#m �c���M@���]P裖��FK����p^4���ٰŗL)[<q�А�E������ q�a��7|gV�)M�C}��B�_En*j��b�a�i�Z\���4�A�g7���@V5�7�_4\�(��S�a[����9���)��;b��·�9�!Ɵ�Q~�C�ߩ#�>�dF����
N ����e]�+�T��ٟ�h���2얚q�κ�����Y�U-�/q\@$��qcE�X�a�u�l�D��^ڤ�Q�;�R��Ԋ��*#���;���4y���? �5���G��.,��_��\p�]?�����/��w(lC�r>f�t_��D�)����5���{'+UD�~����n�*u��� �I�M���m�MV�e��r�/?B.2Q�Ӳ}�x�`��D�Z�P�O#�\�]:�2�DPj<&��sZ~�n�ș�X����o�`�B��av�0��-��`�&a4����f�F�0�� JW���lGd���ny�߼r[�n�c50:Hs7/
�e`Fy�氘ǚ�3*��6�T��ˡT�p����CZ���'��5� Qޓ2VU�FhLn�vxQ�VԽy�Y�l�SR�phC����#
�\�J*�鰠)ɉ�Wф�D�����)����	=�'Ο�����B�_�W�}��Gp�'�Ma���$I��
:f)��O�;�peIk8�R@���/����B����5���E�eX�a�ٜ�Q�n�gf�P�8$���+&ɋݢ�_Y���~�C�_\�̃6��Ƃt�@k��-��ãdiD~�-�~(6'"d�B��L�&,z}�m�4Ǝ���&v�ã#g&��x�T�Od[���jb�bڡ�=� 3�j��)	�������+����q�֦���uj��ٱNm�2�t��N��7�2��V�w��\��y�8�UݐU8!�XEP���{�B%ywf1G��'?!f.���ne��E�7���0n�-�&&Gj��m,ERA����(bC)c@��I!N oz���7�����e������֓՞�?�Ѣ�9����`�?ΠW6�_�b�������3P�e�Kܓ�r��T��͸_�2�y���s#�=b�
Xa�2!]o�P�z�J�Q�֯A�
���W�����B]m4�O��Y���)�\��Á��]�ݺ�h����ShZ~����y[va��gu'�sͺ�KjD�`N�t��2`�w��|�I��F�00�����{/f�	<�V�y���AD�A����sN"��R��i���B�%�����P��ԧ����G�u'�C��Uǫ�L�	E�ݐ�a<�z$�J~A�sՕv\�^�)ῈF@�#���#��*�	 Л��_�����H��㠪%�9"�c%5�è3���A�ˮ۞4�a]ZZ|�r��9Un��4�*���-��f�ڏ�8�n��A�:3M��"�̄���q��Y-�����m���@&R~R!��Y�B=� �Α*q(��,>u�|<E�zۖ�.�����_�;&�h�D}�a!c�"y�sk2?n��HN�I�3qBc�S����CΉ"�	��tif��*,�l}�t�u�I�9�,6� 2ن�R�3X��n2�ז��3L;�b�N��##��3ġ,�zJ�n�/(x�l�,��KB�s��K�Ңq����HDW�cC�J����z�9�<�W<~+9t�)�����,�����,~���"jNnƞ(�$B�p�$�A��˂����tO�a���c!�y��8u�%��s����y6}�s��ggF�~�F��T
�{K�;�7n.э��?�
��2K���տ̹_���F'[V��:Fw�)ҟ(�R&�M��1����,H�H����^��ݺ\��U�疻@C5,P��(�&O�q��������O�����e��F�)Z�r���vj�|}�+��v��k�}�"qʯ�UO3����ٻ�����.��ޝ67}�$-�Ū�H $���҉K<8����N�i�;g�_�1D�p�p�_%�5~���$�CE��*��7<�yLJ�d��ԈEv�t\�k����y,ǺVZ��~�R��K�#!���؏��� 5e�ϴ��Q�u�*��y1 �A���ձ��R)`k7K'[����	['��C���(;�~
��Q���J��5Y�7	������&ꝁ��$��)Nލ�{Fy��o��1���e�Z[[����_}�[3Ҩ����ⷿ{�)�Aeٕ`!��7n��/�	�8I1�h$J�|��~�����S�2>p�ͫ�{�F��ȉ����s�őJqѡ5Jh���.�,i�j�[$k���(�3�����U��`���jɱA�+��KG	n5(���CȖ�m� {��rX������~�T�!�6�����k��<C0�c����O���I����a��ͬ��>�w�5h���봴P�T�!e,8Bi�@+��f����eL������� �����F/�j����Z	�x����ӝ r�{�'QU�p�<<.���
cv�����O��_���r��YH�����$�?Ym�E�L(�s��f��Ĵ[�R�5E}Mk<P�V��\��#�L�l�r��y}�#n����xK���u���k��7�����l�����X�<�1��gh�wq<�vm!�\7����x���&�e$��k�{��l�h�X]1ΝC<�o%Y�a8,a��<ْ�ך�M������$T���Ol�-���c���t��C��V�r�J+=!+������}���?�~�
/�ZF��Q��Y�/±�t��(\�����Q�%#����wǧ�i-#�!�x���}=e�G�~�����h䡧G���eS�Jͽ�̥f����m|�>z�����ڄ�����#���ND��pɲ���Ӊ�#��l�a.����&�DS��209� 3xB�6�4��N��D7��6S��c~�Lu���f6��ܟ�}��~_��3��-R}(����R��-�����ւ��Kx{1�1ڶ����
�~�2˅e�9従�t _��<#H<n*����[���dai�%�iYw�m��Z JC���>;R�
[
Ǜt���.�S�b)�

W���u�a����#V@�֫��_f<0�+ ���։��Z����n�ޔfd��������_a>9M�{����H?�rë@��1Ø��,�L���Gn�+Jbt9S�oh��Y<�0�2;L���۴�9���!��nS�\3���B�dYL�+\��9g��Ο,�J0��p����҈%�gj�f��8�:U*i����V5�}���~��0_��O��Fb��n�4�-0x�����}M�v�lIs�LK���d�( ��k�p��L����e�:���	�vQ�O��*������@?�s�R���z�v��L ����I���|eK��h�Q��&�v�q��k���v^��ޤooG�w,s�1/���bu�������l�KT�5�Q�d��G<�δ���`�B�� 	�MUt��`�M����3jr��.u�%K���V�c��j�E�h^���X|N�¹(u�e�����<7o6�f�G����EdQ��N�,߶\-�R��p(nK��ɟWA�:�k�g|���&��h�X7]��{���5<�!�J��@ ,�Y�}�o���p줺l��4P7[�SXM_�S�$�%eOmas܇��כO���f����^�)�Y�bd�ۤ6f)�����n����_irv)h96$ޤnD��^��+ы��U�$��gk��w�Zȱ���	'��Žh�������U+����$��s�D<I�\�Y����-�H���S�.����>4^��s�@Xx���(:aʚ=#����� f�R[G~�@0En5�6F�E8J���</T^�4Ma���3�%���ٽ���'�O��?j��}����M��܈���G&�ߣv�[�1���)�L#�p�>rQ����H���9�i�c��:�ss�6��B&�)~HA'� `���>;�7@�G��"f?����=�:x)��TR�ZcB�xaBA�7�E�'�7S����S�L�C8���s�xM���PT}C,��J;s�N��F�Q����x��:b�/�y6>n���Nsqr&0L^����/I�w��;TP�� ���@ʣ
��(�3��/�ɉ�};U
�ѽ�v�R�}I����s[�[ؕ[��5|�=�_��I�,��I)g'9;�x�f��)���,�e��Վ�,*�ɀ��W��+U��e�)'x�P:Bp������Z�O��)��0�c�_׾|A��l�nL�]n.�:7\�W`��)j9��#�^��
h�E>��R��eϙ�a�����_!L�oڎ��aT�t�y���(7ո�q��H�&�@��$E� �z[�w~K�0�T�I��G���`r̃��͝S�2e�b�*��RL�96,sa�<:��\w������ˇ��3S� ��uՄ��(��y�
,�p[����T3m�]N/ü���w�(~����u��X����ճ-����y�k������ײ&��9"hn��̯�=�5o뭬�Nl�-��=l�Z70�ƪՖ�Q��Ȧ(� (ҩ��r6��47��OT|�������-@/���]`}��������f�.�����i���Vy.g�>��CQ��*/�J\fU]x�M4�O���c�O��>�g����K4�ծ�vG��,=�3�:}\�W�noJq2�Y�H$�hhA2{���"�+X6D���}���(��Vŭ�y�E�x���^��/q�6�b�Ӈ	�?��I[E��Z+d���\1Y`�7&|�+�W�� °��+����G᱀f"<�hE�V��&�Υ�����l���e���Xg�(�\bڊ"����n��.�k	7O���x�P�}��]4 |�m���^��E��^��L�A�	�F�MAN�Ҩw`,�oi�0m��/�.y���+�r�(x���#�BU,i*���ˆ�LmE���U���2}��y�m�`�C�~ץV�b���o�w��1٥����Tl�D��,�mޫ�L�lx�ژϥh�3�o�fmS�`��� 5;K+]��K��vu����#���j���!z��7)Ƅ�k�(ސ���Ƹ:��{:�#���Oܼ?�:�����e^���jQ��p&�`Q6�J���T�å��Uj%���mw�R�v��R�G^��]	$�+���ʂu����Y�����{�������f��m��o��-��7s��b3�S�A1�:�3��G�#�[[t#M�j�3K�n7�P\�&=�O��T �j�)׽m5И8�2����~H!5�z��	t毯bE��
����w�P�sѱDU�8�M��r���7f����R�)e��No�.-�B<TK���h�'���W&�?7� Bg�ڲ���PQ�T�ξ�'K��۟d&��H���K���qQ]�w��p�Տ���z�XײP����@w�7���6b�=��g��*��բ8��k�,�6-9*yO�*	��S&�EP�!g9	��P���4�MP}Wʷ�b�*��!�3�l�.R]�57�^[ؤ�̍���>��^�7C4w|�#���v�=�aC���h��C�
Bu�m��o�{${��!��F(<Z'�4r�B��}���y=s�6��{5\(����:-oJ��\yJ!i�m�p��������~a�>�Yĺ8���3Z
ʈ�J�z���`��*&צ��b��4�c�	�:�o��} ���=��T(5��rH���W{V��xߩ���;�p�n�h�L�K����f�*�ާS�-c��/Y[�[���E��M��-d3Q_\��aF��"HU�d��p97w�e�ٽ�/�cGwZn���l�B����IaeF	gv��ea��(��2���wش��m�x&u�l���
Dt�] �e�m����`�� �}����ܹ�o^���
C�E?~m��,� #���ͻ�����HV줊�՜G	o����\d1����� ��7��9?Nr<�3�+��`��x~Q�A�l��@c�[�kN���TM��MV���=A�p{�l� 
秚VD�ORH��u&��]��t{�&����i��pQ�V����\�z�}��y�Ū�!U���	�W{�� W��H�i�ީ�W1i;�FD����F]����%�57�g :P��;���u�p`=�E�c|�<�+�<:��Eړ��9��\�,U�W�r+�a�>�-~SBXM_ �ZC��F0�|���`Q�)��#p�ŦKU��1��K�����#�j��M.�3���ag����o$e�@D[m�*&�r�Q�S ����І�lV�ʂ���"�����䫝���r
�����\�;"^H��fc�������8�|�HLƳc��M������BQ�ӗٶz&D����}��$����u��3\�i!C��_=Y�{:
PK��]����Q͛_�ގ{<��J�G6���D3�L��	�kD'����q(�����ߑʹQ��4�@�����\m}RYYs�hT�F��{l%��?���KYY��9ْ�%�1'����:��ăNޏ&��CI��᪾��?g�׺����EX��J��l��f 5V�ފ8�E�	��\���tR_+67�[�+�Gc��B�p�+����P�3a3�D\��Fu�1�6�l(���ᴌ�wc/�t��*�.���ۗ�))\�{�iI��������[>/"$_f���Db��	����d��#"����g%h[G����,P˴�D<HB�����}���%�)�+�LLLbS��m%����2�Ki6�����$k}
 ��`E%ݖ�W�q˾<�=���M�2�P�}�X�C!��������P4�#�b�줎Bd�C$�S�F����hSY�ԝ�3]��V�!�ow��<.�}�[
�� Fֵ���W��6=-/i����>�Wpd��W�X�H�I9��r���	�|�*�mF���]�9�XJjeFE����	�>��2}�,���Έ��tg�#�H���k�����2d(� �C�v��F��`�-�y�]S��M'.�f�����o�c΁x�+`Ywc��#�J��_��=\�N	,�� j�N|�yF�"�o�;�=KH_^u��%�?ι�I�O\֦�e(�TZ��$�zӯ�Y	q�(\y�*��9x�Hl��⣐���A��a��܊��Z̡
m�MF鷾���n��^��r�K>"L��4S<'�d�Q�\�}�ݻ���t8ݰV �����!)������T͐�*MN_B
�!�N2�»�x��Ʒv|��m��eDq>��C4��DE���u��F(�[/Xp�7pօ��Ŗڲ�7j��NL�pƸ���<iR0�D�Vj�`/�Q�@.���m"���`j�ff�G��I%�4��ԍ�$8���X�<��d��7���,NX���Ӱ���)d��q$9�q�O��
�;�A�?��W���!�W	X�B4
�֋^�h7�P=�2��0����h�Im���:VV1�����>�Ih�RQ38�4~^�*A�&(�8�:ݭe�|��a��3����JS.�@%��<E�?��@4��H��OVp���'>bl&�<Y(�����[c'�Jo���p���|{R��2U�5h+Xf,�S
F� �vV�Ĳ�����c���D:�YyY?�t��<��pCo�#�<�^Ⱦy)�9C���~E�����`�G�����5�5���4o>�84Q��������\/Ȟ�0�Q�tQ{���?�W�إ}�~7�H��P?�v�c�zQYr��䛻9�a��mY��x׵�A�O�VF����d"�(5��b��k����^y+��Z)�y���L<�s�rǉ�)|_�T���c�.Q�s:��!�1�BWMzW�����@���2yݵ=��z��B��pIWۛ"�&��\ϕ��K����r�8i�Ɯв��;Z3?� V1�Κ]��ø�9���6�K4�
6�&�f����x�i�
b��h��ɻ�׻�%�;/&b'75�C�-ǍC��R>���_�a�]J��3�FU�(�Yx& ,q+˟_焧D�z��J9ϙ�v�4�;��B�J�zlE����p"V�SI-���M�(���k�W�ea���L��}vo�w����k�����;Z���jz��tN%u�ڕ!{(1���ny���]sy����3^���(�_���00{Q-��!�v����__42�:=Uo���s��O�oQsLJf�XLg*��Ul��\9c,�)yd�_=��9.�������mt��8����7H��j*]i�_P)�͟�q����Iճy�h{.�\����u�/6Z� �N����2�9��l<5{���~��4��)��d�ugb�� ��+�˫���Q����4S��A����_�w���aYz�Iu+�D�dYO�2JT��"Ԕ��Pç�H�9�����츺�s¾H�6�m�OІ��7w�2�)�;�c&
���#V�|�C~���ơ�a�q��٨$HZS@��� ��#��	=��Ɵ�1<bS)Z��Ӂ8�>5�x)��a�Z�X��&���e����j	/5F����d���h��o�D�U@i>�7 >�1����(O6��>PF�y\=JO�"M���I�.�>Z����1,{�r1�F��c]���f�f98Y.���x_�a#^��h���%-Nָ��<-Lυ�� 4R��}�*�KU^�58^��}�g�u���4��3��~�������h\�<�E֦~��9(�^Fj�<8n�fqyu2]+�^vW?��юf��F�:��ܮ{�£���ź�@n�u�1��)�2�0�D��>'�����b<U��嵄�u>��~;��F_~ ����y�E�&�E��E�H�x�����N�8YU-�h�Q�P�:��Z��>=PC�!^�Y�u�o�<�3�x�=?�F��N��0�s�V���XpCyÃ�Wy��;�3��?̘�r��e;�vQ�t�۩��E���F��.��>�S�}[��[ƒ�w����1iA��DC/�+���a%��x��_��(J����h\����(ge}�h� DL�~���r}:�em�ǘ��1��N]����}����l)���a/%�}`�Kg��	�?0؜[Y��k��ȓ#�ޘ�0e��Q�Ƴӏ�g����zy�g9�~�s1q���ׯo|R޺���:�]x���Z�8�^���J�k?��?=D�k�yD��C���=�C���������n�W|o�sK���xЈ�bTlxSp�~_�.�C��HV�p��=��cwgV��U� �_�S��d����}���z�W���R`5'Q��Y�9��9Q��l��r��j3��}��-~���X��^��Űz���F	�}Iq��E���2!Tq�\@�`�=���ߒ��[�]Ɛx���w-�����9�W�X�E�6��e�o�e?����!E����O��)Fv����$R�4>-hܾ=h��N�לtY�aE"ǐ{�a�P(�~�D>���D4�ݰgN ��D(kN��L<����1�I�&����r2�ңD�Zg0?x��8���V�{��Ԭ�AX�r�خr7�A�Y��*׺��"�J�J�G[~�T<k�b�+�M5D�ݝ����I[��@�5H���dbp�B2�8z
��tF�i�����+�H�VO S�����������B7 ��p�ɐU~2���� 9�
��"����x]���"*J8DĶ�l�s򸿌h��o��;���"�r�/��"�����.ɓ]kg�,=��<{ĉ�c���4������-?EW��\�� 6�|q��P�/��j�\��2��st�b���H����.���[�X��l*��o�Pb�G���3=�kk*ܩ������@j��O�cJ���l&I�����Mj��ոߢu/�t�X��M=�%�� ��ب�� ˑX���X��ݬ�����1hjN�>�{����_�z1�]�6%|��@D@�H��[!��=N*�D_ي2�L.�Qm��+��� �_��)^f��I?������=<�$����Ċ
A��_��7J�/�FH��r�(rA؉���긬�0{��
��=G��1TP�Pe�e���?J��o���Եdz�P`B��S��
�6�Q# 9]M�lm���=åA�L���^�{�RBu�je�	��{t�\�q�����(��S������ �/C�,E2��#��
�~�J8��Rt���]2~P;
�Tǿ�����Ēr�ߔ]�ɟG2��Ɓ�%�9�&��g���HHoR���=\$��)Ӧ��K4F�~��'9�@w���}���N�ه���L�B*ֽ���/4�z�Awg�Dz�%{=�sL�w~�:{��eA�-��a��P/G���}��p��w�	��|��0���d}l&M��#�J5|T����rÇ?l[?)Kd��צ���J�̋F9˫5y��K���]�qqȧ��<k�m̧�P=��&f�M  <`Ea�JuysY�Zf��m%6^�@@���T�3�G�M|j|�L�egh#9ӱno�]{�K<C���H+�G��g���pS͑�z����r�e�Bn(.��\Z�5a�2�w��F�*B�	=
�]�Γã����tz��D`JȲ7e�g�N��)��n���\��C�r�H��J1��(��_�TT�
�¡3�/�x Q�?%'*}}
y��Ka�@��5��U�!=�����,B�|���A�J��ځ���zb�1��M�3;v/�A�^9����LV��&����-"��A4(�n*y#����`(:Q�Xp��9�}�j���s�`�T,3�
8˄��������U�ǬՋm+�lYu_YB��*��Hy��a(��H�FȦ9[�<����H ���c(x���F����~~�վ]�����?�60�f��2u�1��ww�������Y.{���1���o��*�3�C�ZLx��"�|y�/�)�2���S
��)�8e�$y��)I����b�'����5�A���.w-�M~���!�����^5I˯_�/3\�+/�.t�=`@r�����������HG��btR���1�HHO�re�H���^#���
���Y��Ա��奙�������~ß(a���?��ՑéPK�ÓD�� cPZ���E��>�Cʰvf
$Ư.�_4��D*g�8d�A~�W�����x|��w�Rk=�L�Ƒq0b8��@��ph	�\@�'2�'<` �%x �\��/���ֹ�vn���}�埘�X;M�UbXx`B�A ���k�׉������������Jx�9�X��J�Ș�]ãd&5z��WtR���L�29c��4|t�^u��Y�5.?�r���tJ�N3�Wn�LY�Y�H52�"���8H�@sT���R1.!"b2��^}
*k5nE8!OM��7��[ ��	-6'	/W�j1�;E �Fs��X��°�����p�S�*x�&nWi�v�6��%�t�:~&���ģǼ
9%�@! �]A����.б�����Ҷ���])���csM�uF���Cc˂�$0�(&>��f��I�8HR��d ����ޤ�Xq��t��1ETh �
-R���/�g�����Ҷ,�J�c�n�¥Υ�ѻ=���v���f?G+[���*�bG|�j�����X�_g�B�L!��q���R�ɂy��>����A���^l�h?��J���U1�j~@���KE.^�_k+`��x��K�4����[Ex��㻦�u�V��v١ZY�ԡ��(����[R�4`wHr=�ex��Z"�`=x��O�X�F%�}��`���~]Ǡ!��vF�Y�M��e� ��45���nT�@��O/��]vn��;B�g<�=�SH��;�����|�%�P$����vp^n��SB� L��,F¤��3�@s*��LG Q�w�x�a��8�e����z�x~����e�"V�r7x>�V~�m�Lay2�MQ�A�4�]`	�1����L*.L��2�S��Ą�:��9�6��,�-R!^�w8t# ���ʸ+�'��Y?�s��0�S"Hk�n�
�z���K��F���4�I�<��!/�0?�Q�Z�^=X�[�}=�^�d�^�1�>���SN�'@���Z���*I����#Vd
c
� ��C��?ݝ�I	2UG+oAdAy�=�U\>r20W�����%>4|�)��7�V��T��[]�i�'O��}�C%�^��s������ܰB�����T ��Us���R���G�`�t��J��2e@\�Z?�����403���Xyq6P�T@���EL��P>������"xϳh�3��uN����č�4䀱$7;�2<͝��n����vH�)��*������C���4�m���ok�������c��r�k9(jЬ/�gUM�&g�F�1�j��G��Mk0X-�2H��K> MG�_ラ�����+i�_�˯� �3yc=��D��J�f�].�pJKj7jM`F�+�����K�O����-u�`֥���$�/�����[��/=�����bT>�}oz�d&K�~��F�s�:,>ʮ@b<5����_C)�tХx����>3H��&���TH�Zo?�ww�n����O!�}�Q�ꄭ�r�h�%h&�~���l�7g4q���o�
��՝�����|� ���SM��W�|J���X��fW���28rK`ϝ��.�����	��?�24����$Q�ԃ{�//��;� �@]	F�'<a���ss�#�kUD7(S6���C����+vbz
á�o�R^��AH��D'qM�I��b���F{?+����'�������7^yPzR�S.:?w�kJ��Jk��_p5�D��wH#��Nh���^ɝ5��,4�d7�G݋�\�>�#�s�_QJpz�TjMb_q>ъ��فY����}�T��,�w��{~�$2>E,o������m�A�mG���)����B��ؕYn!��I��+лd�F>�·Ā�	�];����^f,/>u{%�Fz�)-$��SO�������}iSgLV���ס�b�6ٞ����L�O�i�l��wp���)�b�l��$��OZ��I��ʁ�?�B�y�:����y�jҨ��j*3�s]�?h%6��g�5]0}��KB��JcL���y�B�L&�E�=��^��ůr��|�

�aa����U�c�Q�]Ď���l��)�G���`�G���� �Y8��sv^�8}�0�R�|�=��1:�0�LI����+\Q`٫���T.��B��Jf��ZƓ�؋0{.��얽Ykm�3&7%�՚���j���xd�@Xp>$�A-:
B�OTæ8:�:��v�4Ow�t�f�P����F��$B�|�/5���,A��Q\��\K���_:x@��I���l�����x�/���O���>��viM����*��b+��=���/�ɪ �7�(e%~�r�80���A`���rL#;��Υ��e8Xw�d��҉�Ｌ����9���^�
�Ҳ�뚾m�Յ���Q'��/&>�M1N怸�)�q[���Lt��p �����Ea��&q���{=�\�(���6e��<��W��Y�Ƙ]֣U	�<40i��5,���e9ی��8�Z���.�4��.�y[a�t�	������ӏ�N7V=�������6&%$��J|��iLV*C�k��b!g�؞G祅�e�R��Ң���
̜�
�D���8>��R� ����i4�l		�Mn����_�c��X}��MN(!�3���'��:ޝ���.�\ԫ�_ݜΌ�}��[�
A���h<L���6#~����ARѕ���"��:ƃ�4W�so���hWl@Z�w6�L/s�J���L9��3�<�����&ѻ�;{��֫gv6��˵���$��T|$�S"���<N	���}#�x�l�ݘ�Z�����Hw�Xr�sҝy���4�c珘��� Į_��f#ebgv�V�{T�|�*.��Y������ �üOwG������g�N� q��G,S�b����O�m�&�z��*�@	���Z��#\˽LQo��;R[�ǆk��)��4�܈���:(�2�8#���ӓ-������7�<_D\w��e�tjq��zڅڪy�/�y[��E��������՛�Iʇͽ�uT�g���&�� �r���G���8xL�r�lQ��ipB���ȭ@�ښ�Q�@�����R���X�����oJ�d�������,�e�jϼ�>$-/�ݳ�DpM��qx�(�D��0K[�N�c� �e��s��t�������~�cNO36�lkTZ�eo�[f��BH�?��gQ��U;T��&R�)�<���=',��{.J����&����G���q���j2RׄM�?5��O�d�Ӭ�vF�ò����qD�f��(1-1	p-�^`�~G�*(P��(3r�3*�;���%1����&�9���I���v=R��qh�S���cS���̴��k&U�d��ȇk�g˽���w�A��9y:1��o�5H0�VI�Fݔ��ه}�E�r#V�\�������؃Za1� �Ѯ՚�o����X�I�>�B�\%�=�8��_0).ZMC3k�?M���+=�H�;aP���Da�SfpRP0U�LL�4W02��'Q��M4��f���"ݫ��8uƿ�@��͛RX=�<�|oޠUQ<9��Q;է �0)�.�n�������M�6���*,���t'>_(���p(�E�DGր���Y�f|8�A8��^��� �4bG��p���3��1���~�����^m���24za[dDN����:��H�-��W3w�ז� ��k�37��|>e���ƥ���6�s� ����B�m��~�2	��$�7�#p)$|�]�7����}��a4l�����!E�<f�TG� ��VT�X���xH���G����n���2����B+��$�@�����%߀�u���n��B=�5�,�p�yES!��gU�-�3��{��_#���Uq�)2��Z�����gl���?ӯ
C����U��`N`B���%��q9�.�h���u�kZ�"e��у�zl�8�'�RC{�6���I��]����^�S�$]��I+r���N�B����>\{��D��!?_��e�I�R
lLPh'V<kV�#���2��Q�)�-�v��C��������4�W`8�v=��~95}���l�~��I��Eth���r;���Rm#(����KO�S��[ ���D<�Ԟ�r�����?�X��)��w��Rv-�J���\6+��WWv�7g&�������EB= `���޷y>�ב������r_e�_̋lك��F(Pb̟�k�e�;���'/���ՑM��1���k�{о��OXz(������x�@"q���~"�1z�u|e59���M���:΂�ɱ�I^�7��r��*&�L?��QP\��g)������f#�u�C�0�#��X�����힯SҀ��Qk1Ia�{�S�Ȋ�F�|&�,)�����ΓCj�5�lj�#-F��ˋ��lG(�_�8���BW�~�8�E\"R�v�j#)��}���� �{Z��$����F����0(r���a��o^(�
_�tނ9 ʮ
9�;��]�&�;�j��L�R�E���ҹZ"ʛ�nÚ��vE�ۧͅ�D��4���CeK@.�?9-/�)�q]�ӿ�7�u֛��H�� �'����-�-�e�!�P��Y���	��p�-K{�t�e/���wq��eyUB��L֘��;ޭ%������˭U�J����0i�K^�]��)!O5;��S���K]�Ї�2U��1U�Ђk�&t���_u�tnBQ�-/"�@�x
���!4�H;�15��/7е�4����Ə�N�I��V'�ν�Jt6�w$т&��|��FRw��np�_Mߔ�ěi��,aIhl`����i�l�ڎ����o�|8�lk������	#4F��)��%	�)��+���f(�qX��a4���Rv/��H��͜{��o)�,��	��eF(?�b���%x�EX,W��1Hm]A���&.i����Fo��K���|��K��նU�C���ɲ�+ίx3��6�,�>_߽���Q}߆�}7��AdR���
�"5�L_�5�C�|�[��2���qaz�棜�a�O�]�z��.j3�Yn���ÍIQ\�1��]���Ty����n�*Xk6�.��n�R�Rd^�X'Z䷡�NL�����vm��b7��b�Gn3���RGaSU�;>��9B�@�TVSP��]�.��'S+�H6s��+�6��!Ҳ�N��Fe�c�N=�x��	@�~?:/9&h��5s+M80on߉��E��֪��f]�ެ�a��A��OEv��ј�Z$�5la��d����U�m!{$l4;����:���OF���6�#����e���	����v�R�sf뗞�XS���c��[�V�,O�}$�shn�ӏ��*�����u�9�E��I:3�v5W�K���$��GH���~L�a�L�s��0�,|چ��S[���hg��;�C�`�Y.��s�G݀�m�� �I��c[ٍG��,oh̅��*�zm����ף.TҊ�H��.� Ee�N{k�޲O���<�Ǐ�cOf��v9��cLݷ4)
�j�3����׹�˕��k ]1:�;��߶�M[��$���I��ج)�$����P2N�|@�(n�����Һ�8���E���lڶ��I!��ӆň�a�?�l�V��kM�I�P�Ϙg%n}���!-u%y�Fb�9ȁ�}�Y�����y �¯e D�`8q-��p��򰑋|L�I��n,���Jqz\\'ź[���U�
m�a�s�\E��&�|��E�G��ҷ�Mnt�l�R;�T��OXt`>��l�n�,˩��X�Ʊd��S?xv�U�ʳL�xu����9�&O�y��@���Y(�N��K�Z�?�?ҭ�ǲ�I�(�ya���J������b�P&A��L�n3]�KwB�IՌh/���Ѥȕ�׹ ��������n��(ρ��^������5W�6�S���ֽ(Fau^h
� ���\'�X�y��O�!���aˠDT�N)Q���t%�,f{�s�*,/g��a��zםV���T#���-�UH��u��K���N���#��	8�=�� x��vː8��D�n�p
�x�(�o�
��jg�R�Y�8a,�<���7[��f:�@G)q���ѓh�Gc�3F9�X���\���u�q{��32yo���I^���tCj16V�m&�wr��	h��|ta.3�K��`�;)V�4�]��6���J��&�XT�8� 5,��9�Z����L=�6��� �-&*|4��)�z�6�>��]�B$�9i�
�޹��h���ɇ��yؿ�-`���r��h����pY�6	��H՜p~P�c�\矧p`u��T]Ix=va�#ϵT�
�8���u5�Z́B� �����%�/�t!/{�Z�Ä�wkn�
��;��9�gHzjy<���-U�2�;xLbc��[���3^�x�U��ѕ�@�M�uc��ˬbo�*+�(���g~i�d���(^"�Zn����xeF��	�az��R��Fk``���Dϗ&� �����|c�z���u��k���.'e0ܳt�P��O�^�"%�(�qc�N���Z&%x�0�M����?��a^�PT��(�\R�:��r�s�w�R]$�/�gf�WCE��?Ps]��v���wz�x{��xP`��ŷen�=u� �`����E4��
�"z�(笃�_�����׆�<����?��R�g�sU#�8_�䡮^�_K�U���]�CA0����'�if�8*#�I�1�n����L����.��5�@�3?O%$�G?� ���Ju)/��Њ`��Y�ej���tr��2�z�^YUה��f�NHɤ ٢��.�	}�����(�W?nе�_���>p.�����
�Nm6�`�$�_��K	=Jb7�Ýl��1�k#��o�4I߳t��E�<3{?��Y(!K��\(DU���h�����lybH�z�_��Ɂ�����k��v������0(A�o�h�7so׿q�$v��� ��%Dȍ��@ 4�XC3i��.d#�� K@�5ʻ���
*t���
ȵ�		���_��EXK��ZH�n�%&������J�TYz�x���?v�%*�	�1�I��G��� �/+Q�����?j�!�I]&���p��5�����n.&�/��k�E��Gx8�I�P	��@��,���u��.0$�!��|tF]pt�ΰ�/'�Y���ث��-E���)�# 50xE(X��c��������kG���^��j@pB(ı���JސR�k=�7s��O��<���mUٓ$M _hk�(5$8���ļ��3m�b�{��RM7�2UR�DQ�R���������ޅFH�'�T�g;H��w�=�(c;��^y���*M��:�uu����h�qi�0pѕi�����Y*J�P0�G�?� X�i�c���J�K�<�Q��d��Hx,G���V<|Y�����ǉ��ɡ0�F�C���G;S����r�M�)zwD�Nv�hdd�ʽ'�O��ёR���"����=q"��M�V������������[Y7t5�̥6��}�{�h���}5���D�}�]�,��n`�K:��9�c�Ѡ�e?��Cp
?|x^��_�(���Y�S��f��WgcR��_ �B���c�MD̬G�K��Q� ������
�G�0�z�<�nU�e �$�l�}1�xo��w,�!�r>��պ0�dd7"�gM�fW�(�7�4@{ä�� �W�YR�5�s�K��������l㥁O���TsrI�E�櫹��r�E��0Mfa�04]l�n�������w�?��8f�^��/
A���q8��Dp���p���|��#}Vb�{�8����#& ����"@���܌/!��xJ�G�:�������������̙W@\�&��@�#Ć
�O *�#g��w[�+1��	_��ꈐ,���.����BbǞ��H��>����LT��&ڠ�G�|�i�G�d6�
w��}zy.���$P��(�5{cpV|�!,=�%��6�O�������^�GGfM�ߕ@^��b��~����,K@iR2�쏹�1Q�G���G��y?d'�_Z��jۚaC��%����B�"�p5o���UoL$����[�c}����x�ɧ��x˰�N�������ݛ���)��B�ʓe}a�!�t��j�J�	�{��W��� N����rsOȜ�Fl��r �5�u���Q}�%>3/�ǣ{ ��U�8<����|��gC�\��ӂ�h|�m�J�R�f��6�:&:)}���P�|�, }��k	�8b��Y�+U]�Mq�s�R�9�g�o ��mrz��&XYU��R���5��pڮ=��FjwK��D�u������&���6���~ '-2��(��.y�8�B���#�'�� ,�A`��zu��6N��#��O]n���N�C�%$��S�����K:Mԧq1'�D��Q<�o-�%B���X�n2�v*�����Q�E��6�Q�\	WY�=�W�^����`4b=2�������sh12G!�!��D㮧6��}j�e�zE��>�|�a*�H�ɘ��N�����Ff��Q�k|��k�}��ca��'hz���I-�q=8���L9��NX��&�e��j�(trD��(�3���$8gB��BX#t#�u����b��Mv�:�+m�i�U�C2�K�����ӔpV���kK������V~nn���ħ�����ݼ*t�醗�ˈT��j`��>����C�Q:��	S�2��P��R�¼�~c���1l^���O� �����n��"�a��Q�],��o탛=��d3��3P8��׹1�`Wo��,f���7�+��>ۓs H�����U�e���K̼G`sëF�.�t�GBb���>����em�fH=Θy�W�|�A`�A�G	�ۊ����U)zh4l�5�tI K�lY�Q�ډ�K�m?�Za���EK��rL?O>��P,�$�>��a�hTFװ�I���E�<����q!��+o�"ʛ�{[	�~�)TS�7�3UH�YK�ܴ��� ���i�F�`v��������&}ѣ�X����3�Rzy���@Ŵ���ۃhb��D�&���4��qQnA�fTF�7�'��_H��X%��s=Jw���;	�!&���4�ᘣ�5�Vw�9x=�4�1��䓁�':�觿��c=�/����f�d��ǩ�Go{T��T�D]��>�8)0C���ֿ��J�͊�uW�SD YEi�`(a��W':��6
��@<���ޞ���mT��8�?:����͂��K=�dR,\�5�ץ����.��S�<��#��:A��rk�<vUhA7yU���wWX�����?���f��_����P����̸���W��w��NYjW���Jt\��WB'=��<U>6��q�V�X
��w�gi�jX�]Jua"����;�ZS#��z��#(b&�zSt������լـ������Q�zT�Xɬ���C^I�pSO�.�/�U�y��#L��"ɳ���U�ٮ�(��*�w����'�}�J	p��g\�u���lit�~���'�?�T�<	�����B��K��20�I7�F������1� �y�n����i�����M� ��<zIC*N����E�I,��I�Ξ(�Y�:���si�B���-QY�������d�,L��A$�i.���'�?!�;I '�$��V,���Rp8�ms}?#��+C#��_���^l�&���Q�,�(l��x�ȈE�'	Mŕ�~��*��M�E�<�@8�{��Иս�ǧ��L���;���n�����@��"��t�y��h��� f��q�!���E֍j|>�"8
.w`�w�Q��@�����7��տ�W�?��Bq�๙� ��>A�e���,�-:f��Փ�U�;�	S�c��% h�|Ȍ���'y��OŃG����83������C��Ct�mVg�޸ Q��rR~q��`䬪�2���� ���pI���z�% ]0H�K�/��I"o��Hh� ���CkIr���O ��0&o��yO�t�n\Ǟ��M3b.%{��I�dL \2����v �\��F����2h���]��AsrIo������B��[��* �bI�Y+�|LJ�{>���SN���1/�X��ul�a��T_kM�n\�ִx���p�n�!_�7����-�j�����G����Z�U���=��J�lXϜ@����DC$5�k�ńl��Vj!NP�x9�u��^@&���?��$��,�j
BD��"�I�XB��$�L����Q��ȶ�J���ֿ��7����7�׬�a���3˘�����]��ɪ�D�e���ro����J]����Q񊎌�L��k%c`�s�{B���szySݳ4�?� ��y�e3�K���kLi~o��F#s$�*ݽ+����Wױ3����4�^Qw�#��|�)���k ��5�{�e��v�kĬ ���v�oG`��͙�B��6���+9���9�M챐x��ˍ��8��ǹ��ט=�A��/��-�:�8L�Y���ND�U>�'\�����Gr#�[�z`�=����܃z�����.��bk7 :ݬ˔��4^G	�ekđ@(|]�~WK7���8�;�C�y}��ӝS˫������x0����~y�/4M�vP�ce�^&���M�w�ˢ�n���]�?�P� qN �K� �������xݐޤ������B_.��6��̅I�i`Ȃ�(�1�����G��;hekH��ݩ�~׋�E����ۨˬwo+e)wj5��%/�<e##ű�=�ĺ/��K���nIu5���)4.PD=�@̶�O�	[�3l٘���BdS�Fy����^b5{�[�-��dnA%�Z,`���AJ+|Vp�>%˟V�i��ȆSn���D{�0Q�`z�P���p�r0?N]�jR�|�gq�&�(�nVv�UY�`%�r"�Zm~$j�ƭ��,\ɚ�|��̤�����o	�GS��F�:R�A�SIf�Ax�@c��.;#��q+��le5�C�	A������!/��W>�L8+��!����4��V�D��$��G���E�%��j����w�1�f�ō͛�� כ8�3�&�wk��t�j9�V�.���k#�6o�"q�t:uot�u���F���R�GP��Y��iǘ��x0Q�ڨn���p]����uX̂p��u�rP�� �\`3m�GЩ>XR��N�Kߡ����!+�jؠ�	C�A)α�bZ#h�A ��H����m7���O[�Usk�����oG���������������2p��ZB�CC�����^��S+�2�q賦6�f�1r\�X�M}Qy�nN+64 R�	��]���e��!�{3�h��K=Cӊ&0"f�qq�#Z��Y�WD�PA��ƎnN+=��fI����|��m�ffu�)78��Nakq{)��@2\1g��˃�v�i�rA�8��p�5C�|R܇���3��3�����C����-�ͨ�\2�Ҭ�� 2��ۇ&��n3Q�꠯�?#��i{?39�smX��7qn��<P�\|6l�������OO�2��;M�1�6��n�?�5��l9��//�\�'rL���A �����}�����H�mp�*���T�}��܊0��f�(�����G�T����XU$��(��/	��x��E���d��_�D��u���ktB���,��_>�v��"�6Q��VGi?C��?Tν�SH4�_k1?f�|�ƾ�HH�B��]�75�O��I�\.���Y��s]Fh�X��fc��7�~���v��{��%���p�C�o���5쁃0�u-�2����71��r<�i����?1�¢g��-�*�~M��W%.�נ�"pY��Lk�S���@Y�X�6����!���@������3s�h�9�ٽ�Z��I"����ت�*ֹ�	��hU/���Yypܞ�r !j� /��
x458�3�,���Rqt-"�ֲ��4�!�����u��!p�o��o�T5�j{Rt~���m����(�US�B�ˍ��&�_�/�'S9�\.2n���q[?A�3�W����?CE@^�������'
GM��{ �o_���P�����9�ݫ݃��>$o�m�^9jXQ��Y4�*�X��.O+C�Pз��a�.|6��;����y�nr�2��?yx����ēG�M�z[�l�� "
��e���Z�_ݔ1m�)���J+P��+��`�'H'��pG( ��[z��`�&��"
�T
򸏎E�s�ڋc>O~e�կ�_�6�ms������}��UC>�k��o�D5㓻����Crv��R���φ��"T��-��e�&�Չ6���^��,6��gZNغI�ߋ�\x �6�H�i���$w�mlM����Q�L�n]^15;d��&lJ;���Qcb�@K*ߦKdA���3r�p�D�J����8�c���#��4�Y�qe?�{�e>�o������墖Ї!�*��^�'[m��S����_��X����6f?�G��[=f�&|k�o�Fo�}*�}F�7o��6�0����R�)n��^)�l#w	�|�_�s�ܔ@7ΰ�0<h��(F@��H�M�Q�v{t~c�n�^	����""���lN?��?Z^�j�Qңvm��B��|�_,����۔8wa^`�m{�n%� �7g�M��ўR�����1e�_�΍E�:.k	.�z���yq'�m������lI�
r�q� ��	Ќ����Nݘ��H�NG}������dV���"C����a���\ETL؜0�!'޸��w��y�}���}������6G<���'�`��l��lա�S�!8�U؄�K7���Bĵ�pM��Eueh�7�,"_��h�[M�(�GI� ۣ��K=�o�.f�������6} �g��X0�5��Ͼ���력>��S��0t%�ü��<.�w,��]�i�a���x�)ӆ��f :F#<��[Iș#!�?Q���UU��#�	���~�2b.�G�H� ϯ��}���~�L19 k�b$�,x/�h%!�.;�K��4�k|xx7�C���$�����
V����Χs�9yH�m@ay5[QƩ��Ǯe����D�[D�߈F���>���dc��㽨�q�9?og1w�����[����<-��y&6�[Mb��xB�������d��7%e99��
i�
��%�R�`����ck��S��3�D�<�%0P��5���UkϚD�h�������Q4v�zψ�2���������V]\E��9J����n��P�l��+:`�[#���3�["���x���_���:h�BL�HM����}{�Q�����q���=E�ݳ��>~�K�?�����R�<�N 3���&���R�
Pɍ����E1��^�!l���s`�"�#0d5�<<��%�����i�& +�bH�p����p���W�B����	�u�����j~�{�e�^�H){���8f�P�A���M1��])��4���sq1S��ȴ�o��d��n'ƇJ�A��NА�i�j�����B�8�������ܴђ�j*�4��(��u��%�8��2$�����>�E�9윗l����荀ռ%�+n���p��~^��/� ��}B�[X�Do�4{_�pb�HΦ�����%L��W^L�j� �ܢ��������=!��۩����ۭ�ϸ�f��k5�Ws�WB�{� �on�g~�Y��W�������%�:EZ_2��}r.�Н���\d�������5���C��8Z����i��:�P+�<�Н�gp�JN6V-N�x�ê�[���ԃ�1���[h���<!��<�f\'&�g�����Bl��\��صn.��SniH[���~���ɢ���.��y����M�Z�L�
��{��lwƫ�_7�E������|�j
�Z�b�i��������э��hb���
�"��i�Z^t�����V(�w�|�$f3���Y�cMV�����U"- ��|x����%E՜��H$�l'��,1�8f�t���Je�*�O(�S�ǄJ��v���Y��bWz�-�?_�6�et��/Ez4n)fӐ(�%}���E��P��ܫ�D̯±��Eh)Sw�q���ؙV�Q����wm`>�4�f��*{L_I+ΰ�9s��-l�f��x�n�s/I�Xa&oN��ױP� m�$/IZ`q�c�`1��c�!�����+�kz'k�K��^�����]W�_Bl� ��h���Ϛ��J���x���g!e���,}`�x ���\��E��&L~���EV��ִ�1D��b�������j��5����c�Ak��{i�eT|�[44�r��c�����,/F��M]��	=_
-��D�����T%G��_M��Rmq�_�>v�$�2�e?H� yo#�8�3� i� YD&)���V�H^�m�<j�!9_	<� ���Y
I���ٺ��GQ/Qm��oXQF����g@�"�����Cc�ܣ���[���N�>� B��~�@��ZQyԆ��QZ����p &���`S�we��ʋ`y�Jx��-�U�^�3$�Us��z�S��Ëm���/�o�*���W�h?9�������4?>7��q�v_@�KT�d/�f��dǝJ'=qy"�$�'o����j)�ci^ 螔�U6�+*�#2�{}��z�����3�^���J�-28��v�_��Bn���t�y0�̈ݗ?<�9b��-QN��n���M �d����G�����H é�����7��HLo-H�7<���c������h��W���RB�<f~�1Ye�C���Rm��������w�E��cuL/X�/rr3�ý�׸%d#�%��`&�	>hiI��,��:�`�-�҄0�Y��;��\�i�Oɽ�To�b�Aɛ�����l�)�z>�
��:���),B��'�fp�2`�,���T����p����B:?7G��E��,��y�A����a��Z�����|��2=o�T�K���xB����a������6$�_q����3�!��1�a}��W��d�3�T�3�_<~���Rv�\��aTLSj�������z�u.&5H��L�
�N&|�n�\7�r����sh�D7�Tèճ�5�؎w���)��	 #4�1�etƣ��J����a�5�����Wc5os����S�%6�~�Q��l��p����i�GP
��EV��W��
%��l��Ji���z{�_=	�M*��:E������1fФ='�j� �����՘�>fp;� \b��{���WIե�&�t�־jҔ����0z�XG�0��a4��3�"<��m`�ls��7V�EF&���@�IN!0��6�t�Jթ�'��Ӥb���H�	���'��~��P��o!���b���r�I1$y۲a6=��v6��|	�ȏ�9G�����@�Q'bW^V� K�,lƣ�ڮ%�;̷i]�����d�9��֌L����T�����2�����1�\)�Lu�1�j�Wٟ�I�U[YOm�!m�����Q��N�Ø����?RZM���M�R� �J��}.ܓ��#�����2�)�,陼�e8��c,0/$_�M�e�(!�����s�(�ȼW��6��0߁�}��Al�e�a�;m �"���j��,o�z������#%�)�ש=}�sq�7Ί!kܬ�p5�c��b��s�~7��<X1'�5W�	��/m�r�b��GWOWH�C;v�`��+����S����O�F?g��q�ԋE!º����	����c5����A�T:C����J,h!t-�a@~J�lqA��Me@�ňգF���r�y$�Ӽ[Y�s����hȠIe�xN &��H䭤Ij�~�bJs�/�CM_\����y�ؐC���4�ݔ�#��R�Ƥ "au%��_�l�6T=�M��0��a��ˀ֢�RK�*�B��J����_'L�+���7ٔZl� 9��c3�Z���B�o8�ɩ�á�^����mRŉ��%��A�;{�@��Ꮕb��]q�<�a����J�o������26��WB� G^8�M�Yp,-�]�.(��Z��)13�<zi�8��It�=���3�0�F�Ѡ��vϡK��5����pWd���H��o���ih�3��MEO"���B��FW�`蟣e@Ȫ�B��H��q_瓄�d�(�&~��oz��6��������c�y3P�(ŕz�lk�i���Ա]�!)6�u���Sմ��H҇^�*� �{�ľ�i_@�mu_�]2�J������<�h����"�{L��6J���}f��
ۈ�Ȗ~.j_G�&r*u,�/���M}�e��p��>�����F��=��Qq�
���rU�$�E�Bz�ѫ�kkbZ^ƶ��i%5ű�m�}��9]GP��@c����(�s)G ;&�K�W������j��fz�t��O�Q�#�皟@D�\��=ٓ���g��~2��Ԭ����o�ư-����/�3($�A�C�����Acv�%���ά)�x�ȞY8#�W 5s��+Ux����u�լ�Ϝ�x�� \[��if�� D�|�j��U&R�a"]�u�����,˺WW$���חWi�kR�h��Ex%��fܴ��E���E<z�#O��3��t=&6:ϧw�~�Dtx�rx���"��(��U흄������g,e�w�ݧQRyf�j�Yl��p�lWm��)ZE�@b$Q[�7�#���
Y,_Bf�4�TG����6VL��������j�˘+{5ګ/1٫���Ȼ�O3�x�ѩ���:�zv�f�P�����Ѧ�y
��W����a���:�u�+MЈr��r�[U�p|.��O��WYK(}zk�UY����6o����V%PI��( B*�|{���c'-��-y��3�^/��Qt��1�#�90pu���1�<`�5g�>Su�%��i�xI�Bv"�Pw�5�' �A�֔�����#6ܑ�c1�9�2oM ��5��R�y��,ś?�ێgӔ��	d���{��S�w	L�藞c���Y��`�ނup�L�����Z�N�Ak�k=�]?^�N6:a{� h�'S�b7���\�%r{�RV�sB�� 3�]ϔX����>�����`�h�K�0|﫫�W'~,�����.���=���̺�/�x�";�`=M�.I�"�
��7�(��/�ED=��Z�Q>����Q�����V�+��/jq���e{9�]fX�<���bsUYbb�G��^c?�<t�Aa{�$b�]�.J`M���n+��?��*R"�EwwR�yF�@��3{ލ�U7��Ť�7{N,�2o�:S�o�j--j�v>�e=ג��-F�hi.H^�q��$�\��tR��$`�yqM��ۺj��@:��ɸ���#��L�ɜ������V"�1nYRlo����u�>�R\q�P�v�Q����/�
�^��-�֛���H
�!�D<yi�)���9r��z"+aƟ�$zA�t-gJ�<<Wco}�66*F�ǉ���be������t�Ǎ��d_n��"�Zb�'T����I��w��v��QgCn\l�(���ӻ�M���K�|?/e h�ec�섾�b�b6F���f��у���p��oO;.1%�7c�H����1���^� ћ�{4�$�3���{y��x�ہ�� f[�����uH*����#Rٙ�����$>̩������z�������	g�h+�S� ����^��_�=�
�6��.k��j���u���'��^�㺑M��螩����6p#l������XE/�>M�Vb=(��}m=�a~�Ex��E�0�ʤon��+�=����q��}7hσ ̋$	�,
?����k��rI~�z���$&@�|ヴ��Kj�`�D}7<�J�j)�a\���M��כ��_��n�Xw�z
�PUȐt>�0l�q��V!]���nQ�0����nhR���F�&�!9�s
�/�������1Mt��"GNr���0��)�!oh��ۏ���j�U���v�V��)NB��Ǵ�8��ח�Ί +��N�.�a��"U��*��4��=��MC�)�<u��Ů-ҋ��C��;4 T��O�B��%@ZvR�c������J��� �>py>�w���Ay����kvc�~���	B��~|�߼��2�vĪ%'X)j�=Uϗ�26s��?�$
lou�(^��w�c<��V&�AC�B���R�6%�x�����YT��vwD���F�Z�5�4����0'�Hꇱ��Hb�S/����Z���\�[^k~s���卑<��Ē2��	:��U	�2��� �/��_�7��񭽮�� �D<'_�����`��\m,��m�^A��3����!�K�薴���C��N�B�Q��� @fL�CاةA��Çx����]�X�о����d�:il��;1�T���
�=:��P4 ������}A��G��hy#XA�.,�
�/xc�`�_�1�L
AK��~h�k+٦�z居��q���oUY�QB.�ϼ�7�i��yQ�I6Ŕ�B��������'��J���h����f�>	�I�ESx�q���m�����XP(A=��g+�Rh��	���KO��߇�v���1Z�o����8����va�\/�j`9�V�3��G#z������|/?��A�<+$؛8@1q>�+LR(�ud���3�J��AF�� ���~D5	�Xs,#�!���9/�%2�#(��
�h�[�ю��8n�wW��q���Sf�?�B��]�r�0�H��h��O}H��D>���2J��T5x�n*��P-1��:�_y�Zkf��ty~ɮ�oi���q}��E<��B�D�G��1� �P�{��x_'�~1����dC!�c��ƚ�7�;Jj闐�����t�C-s�Ab��0� WgDl�c�_?e��Ŧ��Y˪w��:� ��c�u��	�QkwO�X,uV��~
���lR�����h��5�Ik
���+d�OHFi�8;m�qw���>�w���gN}s����y���q���N9�����������D�l?_�; �55�4hR���kI3m~�: ���[�bE�m?�i2θ	��/�.�q�gH�$���
�?qI��C OF�Z��m�[۝$J��q�_Q�ͩ�\��?�G���J'J
����Y�E�ƌ1��Ϗ��[{��r�1�T"\�����35���)fPb�����O� MQsPj��D6�c6P����:)ץ�a��"�K�Ng�+tVq�YY��kB��R��
4�Q�a�ii���k[H����Wb��phX�F�>�lI���9�YR�f�`�h�K;�_.�yO�N�C��kG���k�Tc=��Z2�Z����d$zpp���[�a�_���	4�ǋ~Q|�vOB�U�cr�/�Z�
^�trԛd5�t�'!���`'i�S�)S����S���� �������',\��t�ޝ�Щ���h�dD�Ax�����<�� ��06�J<���Byy}-[��a��2�9o�؏�*ܸ;O7��U���B�H:4��|t���!�nߨc�%*�POaQ���G���p1^���ٖ�mq��Tm���i֭� �1)_d�鮵���Lt��}E�K�4乲���ә)�&ȇ�����o��b|����5/׫ �-b��f���נ��!2�� �X�b��!y�(`3��=�GU_>/$~�/���`M8#����J�P�D���'��d)Vl?n��`O/�����(�Vj�����?p]���J %��:�`{�?��[�TJ�	o�	Fk3M� ��O�b��A�-���S��k���ǡ�ʲO/�=�
#�R݂�z�l�w{��.'��Wb��x:�M�/g��k��3/��3u�������A���A�A��}��4#y��j��O��:��_̘����v3`�ը�#cÍ9='��l%��� ��;��ޙN]`�]��Tj��1Q�" ���E�p!-�*�w�T_��]V�U2Z_��,����N+h�v�^��C���\�����^��m�׆���¹JGT٠$\Gn��4�JM�S3i`	V��u$�ros��trʄ	��2���<|uv7'*	AP;F M��*8$��ŴO)i�VH`���A[������6��I3T�.���E���	O:�x1w�����G(#�I���2ˇ͕�e��Ʊ��ͯ,�9��uс��HYԁL�	�@˩Mdt����/ .�ؿ����)`0��7r��%ᯛ�S���ޫ������洰��vFn�l\��]��^�cn����!�(/��aJ�u����k�m��C�M9��&:m��=s��bR��?پ0%A^��A�!�R���*KA��e8R�*��N皆�P�iDi��1�z��w��H_J�4�~�58@�\��P<T����F����u�v�*��d��v�+��#�s�F�_zH���ڮFb��iP��w���q�s{��[I__:[�/]e4�|�W�)��d)K����T��V`��ɿ4�5�yHN�{V-w)���µ%
&S�������4Q��U�1&�ӧ�9b<020]���K�5�|!fw��<���x�a՞���H�瑲��".��!:k��'C|΀���P�=22n���J���V.�uA���wʪ�W�Ō���UCA�a��S��������4�6�'~S<y��E}S`G���T]J.���,+�uU1&V;�$�ت��[�Z:$
?M5�bSX��[[&ׅr��$�.��nZ��ԅ����pV_{SPSoD�zV�й*��;<-��\����⸓8�9*J�:p��t��h��Hm�w��݅�ٵј?̾9~�Gx���!ǧ��)����g�8V�-:ͮ�+г��`C�6-��u���l�%�����`��;V^7k��2a��Fb��!�&��:2`3�lJ�%oy�=�������aR��m�Up�i?)8q�`�I��m1�$�Yb��ʠn��S�K��J5[�U����C�ճ��[d�c�K���jW�cʱ�WVcdqoq
W[�@��tڙ;��|������/���x;�o�,3�Bp�N:��0X��W��S�H�r�[`۹����5�`�௑B���M�^O�ZU�Ԙt&�Aٚ��0�'�-�^Ć}}�(7��%��c|FD�Y�6�s:9��n��N���#H��1f6/x<�2vKW�W����R�<�%�ޘ� ��8�/�E��1ic4�ȑ�:� ��Y��:�c��"rү5�{1��?Mτ����"|�u�B��F�)�TB�5
+�_\��38��Ҡ��Z�.�~M��K�s��h�0�$f�ե�t}�����]������"��B���ز��8��ʬ;mwTE(;�`{l�m�������N1i�/�R4<�[р��1M����4ZZh��v�+}�?���fn�d��30���`
��0d
y��RmOqw����MG��Ӵb�~c�M��#���^�ښܨl��^�l�gO<���g��	'F	<gV�{��@��n�����sY�z2Q�*��pXsK�[3wm�\o�d�HAF Wq56x��k7B
�~5�����Om��q�*�@�� +g�ʹ �A�c@gm��+q'sA^����v�����RP�ű�e��M���%wp�	iO�ol���K����>�(L�-�����q��`��f��`����˛�� �D0�f�(��)�omd�긖������Lk:���A�"�F���#�Ji�0�>��P?��Uww�v&�Ή����a5��4��ʀJ� �\G��:\��]-^�t���ݾk��N5 �9�3��f_�C���4}Ԭ��`�y�|e#���|g�0N&�x�1�`͠�@�G4o��p�s����ϙm�+��т�Ojb� �@Nk�f*��N#t�����<w8څ�ek��c���� ��冸�Sek�V@��)BX�aB��=�� �ŝ��R��Ŕm̜�ԗ��X�̗=ʻJ-�?��ϰ�Vw�>
�a22Q�w�<3�A��'���e��i"��QT�K��f-!g[T�l,x֑^٪'I�K)���J�@�4V� .�mG}V�7 &˝����(xwΜ�������������'4#}�#�/*�Ak��s+����f�Ԫ���,���^Z�U�@>}b�3��\��?�E�	��Pʣ���<���@q;���.Y�>V�.�qM�ц�)�`����i�X������\�+p���|�+M�oGb$�k�^�o��L��=�M�@Xzw��L=��5�k`���q!��Q�k��	>~��=Y!����w�D�|B���>���\�m�#�̣���;�h6[��%�
�,<d�g����q{�jY�%��W�cЬd�/�v���=��O׹"ra%�y�򀓵M�F.���u���V�M�j���~A���YL ud���[���U5�+$��=���f;��Q1$q����q�ȑ�6I#h2���y�{�:�{�r�ڳ�k��S��_�����Y���v�����R���\��)�<���L�T������$ߓO��R,G��Y�RQq.n���ܦB�=�@S�� �]���S����{?˸�u��m�U��Y�8�0�
��!�Q��'��k���p��n��E�D�X7s){�(R#�*#�M­�?���3�W5�秕�^22�}�#}ҙ[�+���v�*��t:�V�Q��1������M�`G_��j[�	�^A?�����'8�㥱KV��r�Q32���,룭�>u��?~�p%Z��t�&�y�s�f���\��3��������3Uo��v-��h2([��B�
��ڴo����t��u�����ב� :�����e ��;]��HjZ�܎�P����oن������X�PZN�$��H�=�5��c���,��~�SS����f2�>k.;j}�t���Rf��ԲZ�e���8EA<C�[�]�{a���/��	x|��i�+̜�rUċ�r(���vy���oؒl��&��9mQ����M���}15l7
����/���Z1�(*Ԙ@&�w?O,�>�$��X�NGئ�/n"�F��l����_��}	��
��LbVl�饽>q-q,����64������\z[�B[ �4 ��2�y
c(wbjn�&��e�{z�]|��s]�; ��:NPҾ�A��S�5�OD+_��I�����VV���M�a����%wn�����QOf�TO����)k
4׫�t�5�N�zwrѯ�v'u+i%���32=�^Z8%�W�-�I)s���t>�"��k�Q2�f���s6���]W�H���GO�C��\���e��`���v0�*캞N
ٰ���{",�C�}��Y�Cp��c͓x�좻�u���Y�6�� ����dq?�����̠�ǔQk��q�1B��"���E]P���h�����z� ���#f��=�'H��Ff���dB��`�N��mD.��_hT6~�:�핟(\Z��i�ئ�{��\P�i;��E(�o�����H�8L%�z�$,x�h��d�F�����A�\M��L����ޅH��r��Q�`��wi��h�U9�aRi��x�T[,^Ǧ.	g�����;�*M^�H$|q��*ܥ��O����n#&�oڴq��3����#:�vһ*1����ck��՘�Utk�*���ȋ��,�ާ�ٝ�_��#�}|��>�#��~��ezO�Ј�٦���S����m���UP[�����5���:P�ؾ6}^W|\�Z��b���Ze��i�TC$��g:�e2�DeQ�0�f����s��M�[_F�7g
;̜c��M�.�����J�rc\<���LG�	pR.�W�e�q�!y���$�C�v�^}�$E5ȼh�ɗK�,oe(Qn���,�KCO��"��ޘ:�`� �������@��3G1H������o�4siK�����R����x~�Zg4�@ssU���fR$9�_���͊�R5������<�é�C1.�8�<�Zm�g�P�����J�]?�&5�"�N���,-ygYEPf�y^�5u�2����&������JK���3�Ѡgj����ް�|n�-��Мޘ�Oh�����݊�����]�
W�J�!�V��;o��g�aF����K���=c��x�ÍH�R����4�����!&Dmj��`q���h�Y��Q&�v{�*缾.vWh�3<�g��']*��aws��^%π���:Ǒ��u������B:>}��r�*�4�k�t�R(X�z��^��֡z���t�,�o8��Ez�:n�#Lvg �`����]����=LY��	��Q��^�����x`AQ0U)_e~��7y9��9�����5���X�s�e�����q��l��Wt��!�!]��X�%��#��Hv̓վ����0�P�$?u^J�����!�M��=6�Q��~^(h\\���Er;дP�Z���ƾ�v�IR�J���=ڼ&���a�BEo�l�]x�|��h��N��Q����SA��{�}����ZvЛ�ڇa��3�z�g
>�٨2�z�����3X��V� �׭��ݶ�5�9{#���fB�~�鸫�2f���,��v��]���td8�7����>�5�k���j�p��2�Jՠ�dL�h�e�!W�r�r�X0|�L����]�����y�������+��=K��U:����K���e�Y�vn�*��ؼ;��]����3��A,��)N1���k-�C{���*�a�AB/pф������3ݜ�qY�|������7+R���eQ}��׆�<1�(}�値!�������J��,� j{kԿ�`]�ԕ��S�c&��U�{pt\�ґ0��ꓷ[Y�$�������; �������]ī�e�Cg�>W��L�k�r�c6c�l�,�d�?��jU �S�g>��e��=�M�k�3qwV31.;7BM��)�t=��&|�ʃ	�����j���> �� ��#�sB-���޶�F]�*�!~���ބ@梡�*`���Ԅ�dΪ�lq�L�*��$�%��_o�׳�<��1(�B���k)x�S�ͪ��b=#>sF �t1~��>n��k�H����F�HE�,�~�46�u�xb"�^����Z�*�p�V���S���惿F��oD�Ͱ�V�X�^��07��\�@��N��e!���S����$�µ�'v����ݡ��X � � F���R1�w��)��\/v!aB&��RWi��'�HG���W��$�� ��|9��Rh��dGN�}MVE8�kRPr�l�7��h��K�~�ά�*���{�:�)�_$����o ������3��1;�oMI*�n~�u�>�T{ȴ-M����>f����Ɛ뀉��̏��C��1Z��~���i.ΐw?�8,Ux�@0�EIFj�Gm��e
�o��Y��E3���܆X�&��e~����I���x�2�q&���jF爪c��Ewy�4���ۖ�^>D���I�[?4��,�iGb����^L��*ȓ�l�jr.�����PE����_�����i�fsMB�%�݊QP���&��������Ktv3
k��_wz9��?�2����k��"���S�^�]��PJ�[pE�>�����܅��>\4��A <S��[J��Dd8�4NU�ʶmH喩�+*�ӷ����Q�{�K����'�mY.Λ�ߕ���'���0�sT�g�oa��$���b�Ӏ��K��;���ͦ�1�М��?Z���>@��<p$�,���%R�M���*u�����[���G��K6��ݘ���2�\������B�&x�Y�pn�$
�xh����4,lI9ex�T�yں�P��J/���tą3y ����\�m�3H�E�G &�����P^����ؖ�l��s6��x����r�]��� l�,CH k�:�z�;䫺���K�u�3��㹚�K�"�bͭB�����z@�0eQ��*�о�W��[6�V�z�z��z�Y����@�'lT�ן���7#F�@w��e� ����zTcl� �}Z=~C��b�@W���z�g%��]"/���&�r�(,?�9|����#�_S��@�r��3��G�5�$�>��U9ί@sv�h'�Yu)n��"����� Rǘb�9 5 ����A�G��$E:�D�}�I^��4��%�!	7K5~S)x_a�:<3k����L��;������1��}����UA�o5R��/�&vgX�E0�mZO�0E��ս��i�7��z��I�}9��;�:O��ޱ� ظQ�ؘ�S)��]U"�k�	��*��5A�4v�⷗��_�(Q���@
�{aU��m���ɡ��{a��&Y��ؕ�ԺFB�1H#��殽�5���b�?.KV E�g�3AE�ͷ�����q���Dɩ�����G�U޻	4��e�J�Nc#/�P��]V�"��K�2E$1�+52����"�hs7�9G_����Yļ����0��3i�OO ���d�;�R�NR�E�YaN$��f�ҧ�?a�xo�vxJBZ��柛��|.MY9��ٕ�,��K�U/�2��������F�O�M�g��E��x]��?<�p8(-f��mP#`���Y#�ڞU���k���;����7ɲ\�J�<���M��@F��Z&��'�A�αl��ޞ�}�)&��i�+�yӍ�]����e(7�Q�90�N�/R��M\��M���0ǡV',X��5���>y�D��<E�
W^��Ո>�����˗���^;P�*N�9X�>o���S��TB4�A-�^7��C��d���nh����SL�G� }{�}�UӰm:��"r2���M��,�A���L�Kݺ��h0�}�\��4#���/d^��լkF�[�6��	?@c���2��h��V����G8 b�J�?�T��.
Mn�o^1��Z�6���%>$a*]��Y��> *K�"=h�,S.�;r�� ��M����AAh��?)�6%ޣm��_-��(^�������GF���z�_��٬�t��$��^��a�{%���yt�q��5yq$ٟϋ����x�[;�DI��2��E��*��&@d��#l#'X�LI�:~������$4�d�V{g@��I_�������ND��H��#��w��=`dL��I{�����o��͘���:��bS/8�B�q߾����B��u�e=��9߼�j!\;�@b��D!�=($I��@�RWgU���s �����nfq�e#z*�Įwk��1�����@�����<�a6QOgz��l�yP�L�Df�YK���m�m;j��q>���?�����wz�˲�2؏[]�p͡�@ϓ�*��Qڗ�@!H��SG���Ɛ\��<�a.T5d�w.&,�/��4����H��Q �F����X����Y�O,���"2M\G3 �KΑL ��e���;��߈��;�sk\k.��>C�g��sy���r1RYW �Ј�����]:��I6A��%r��$����$:̑�9{p���hYޔ^��	fҐ�OݳW|�i��ZsYLAMC�WP�j�s, =DE-�=9�Ɠ��| 5�[@�q)���|����|S�f��}U�R�b�&��'����۬�!�U�=���%���>5u�a>�R����� D4�=܍��s�E',����LQ�c��p=�\C����-Y��F)x�/����Q��9�(��$WH~�}�QÍ͈d�7�o�U�����1�Q ��S�wwkp�G;�ѐco�̘5K�WB�����;D�/?�^4BlT��no�#�~-�,i��A��GM��2"���E��<]枎Qe a�E�b��^Շ��t+7������w�~��*����R)�����n��� ��;� ���~t*���b��aT����͒���M�b�����|;!��#�Q���զ'�%���}�������5��9�O���<n�Q�d�+���C�Q�ΝoN�Bɛx����Gi���ms�pPW�����nI
d���4C��wg�@����j�id�0�o��+����L4�i�g@��!>]�S�$^;��3���>��P~���Il�,��l������B>�R~rem�H����`{E�>��}��+����}��aXӫ�<�p�[��rAOf���/�(f�z!�j�����Y�b�r�>����	�(�4�T5���9Y������W#EMQl�CTA\mwg���o`ꉯ7K�-=ge��O��L��>��[��=�/�[4���4�0 {����m�Ѻ�|s�Tcg�{=�ɠa$�,+(�(��~����S�Q�=uQN7|6&*g���X�a��ky��u|�<Ͼ���8�J�)+�-I�:��Ҹ|�DV$pjD@	;����o@[�"a[�y;�)QT޺z�v���Z���y� �:�Q5
���;�z2
��|���'\XtҊ�N0�8��zJ�
�*�?h���X��^¶o>bch�9h�SD��	���������M���Y����-M-�]��a���G���+mN$s�h)��"�^`z����]!Ҥ������P��f�l~4��3��V�& �S������*�����D>�*d(��	�!��{���l�cv�M��c��sOؕF�R�q>Rb� 6���%ơP.�����R{�S��߽1�7�yPQ��);Y$�Y��k:uČ��e!KN���U�KÀ3Cr�i?�W�ϴ���b�!�u��Yf�{��蜿i'�m+��]�Jv�*W��-_��/@o)��Ҭ����tߦ�E3�������|@<t<�^��PC�^�]��^*�N�FA�&M���{�]G���d8Q�m����4V>�*c��� �!�o�-�3㠂����y��]�&�R�VJ�Ġ峀<�B�+E�WG7�:�S�	M�o9���p�[g��˹��z-fuS���)�eb�������0s�()����Z�D�i���m��E�)3<N�r��؂�Rb��զB��D� 	W���e�+�%<���c��6�.,����+%閩�O��sP��4��]L�h�����;��LA�]�2��{����"�^�5.�0j�[Yӈ�-<u��)`x��O<EǛ�y�si�Me��x=�I0�:��`���C��c�X:�Hߐ�2�r���q�ǛǊ����Xse�w�������gZo6]��{Gbd�AK�)�IW�Z�!���<�w�}0�hI���2"-X� @ �<ֵ����[�QQ�n�>��s��3�tm�B�,��_�ק����늠&YK���0�;��#|�u4Ѵ��xԏ�1;9X�h��(�f.�M��k}�ߵ>ZJR���!�Ք��[��#]}��Z�!��FP�*���<~)��S�xX9�ۙ�G�� �T��$|�.��)�s<-�6��ؽl|�c>�PTZ�=��/������v�6�eUz�����T�������!7�1*g(�]�.�P ّ#α�A�Σ����;r�g�v�v"F|�ז~1� �T�Wè;�ς)�&$�
%�l ؞k'13�Q��윃?�fQ'}��>��6#��$o�z��0�RͦG��Jq8�!F��ʐ�2�ʄA�Oh���v��*a�Z�������@o��7���y.TsZd��w�y����"�&���Bg��Nb��S���Q	ՙQ���o��]C��WR�����*��4Uy*���ƨ4�;�_XCn�\C��,ockt�yo���V�[��Ӌ����������l���h�9*�~'@K��3dU�&�]"wm�(J�j�N���瘴�Y��Ep�~\�V"�5�S��n��O���zาm0(���Oos�z8qTܼ�Gt��Kc�Ӡ���p������p&�0|q˧�	Y�gf�P���*wΌ�TA�&��_�8�^��������s�L� W,H���Y�p������m����,ސm)f�\��U��1�O��}:�:<O{�t�zE���N}?R+�A��ߏ��B��yY;'h��g00����X�sI{�)�PBΒ��p'��L�]�f]i���>;������p�Z�M^�+tGI�h���
�2EA�+wSW�K�R+��ۗDuf`]����t �mѸ[4�����j�=c�!Qi��;���Y5E�9ܶNB��ÛG��Φ7�H�-=�����y] �ӵB�dr�f3N2)�'ቴ�e�A���+?~Ձ9lK`��U8 VU֥$�B<e��]���;Kҁc�)���G~����i��r�>��Cܗ�3�.��{E�x����q>�\��O��zv���͡�<�ω0F����f��qۘ}AB�u�&$C��x��IZ�`sXM���2W �Q�mW茼;b�4y�U��a3�����b�e�O	�c.�Q��Ihc��X��8����ApW��)���2Q��,���_�%��[�I�����.�fupT��L� #P�:62�'����4�o��S��lO�(wx�E�.�^8MX�o H�������"����W���^Q��1��L�[�]�L*���y9���v3=+n��5��=&=��������P�e����߯$������[�g�8�R����Hn-=����v��U-sL5~'T�YXqF_�+�ASc�Kj� �GA��6�,F"���������r.a�['� �(ʋ�%����ٽ'?�xR�ي�TeH��d%�/�<A4�aǑ��C���U�']�!6��o��1G�:CAjm/T� iXY�d����*h�t��g�Q���{񯟣�u+ܛd3���������nX��N`�� �V�`�u�fjT�)����x/��+�p}�zO�PߝH�J�ޏj}h��Gnco�%g�u�e���F���hj��8X���+Z�_���W�{'������s!)Ⱉ�����"�r��x�$��B0�S���h�Y��(vc���c{����#ƙD�X�A��}W��9����E�78xY�H��(#�õ�]>�=a�p��>�%r�]M��H�o-�'/��U�J��ɒ�osT.8I�X�O��M��'���?����g��������33@���}]<q̉�I|�/I�N�$��CL�U�R�JB;ur��t��+�t�Cg�Z#xR�9t1
��ğmiå�bw�`E�eZ���8��M�	��)g����h�ΐt�44w�r�<_���������n��u�GE�'p�Y��a0����<�"3��8O~�e�jn�g����r�up.�B����A���,>Ӵ!
͐�i}��t:�|�oE�TNW��m��\>٠�F�H��?��N#�N��휖�V<�wXЂ���P������73��)����W����X{��J�xB�4�����pk�UX�dL�f��Z"-�G��TQ���,�(+�R��E�*��񀪒%�k�D�����;^�X�
���14�QKuoNC�g���K|�G�*�}�7Bhꠠ7�w���"���02�]K�h&�����P����7�PĜ���j>��uHM"�7�5\_���:�02��M
Y�-j�$�)
�/�$�#�2E}m�UQ�w�c�n�D���`��Ot���Ԙ;N��)�\�u�ܒ���S�Ќ��c�6����P#Ҡ��ɚw����Lݹ�^�4�<!(�s�j��/�H�D�5�IJ���޹�c�?^"��k�e�� ȧpF�d�׍�y��c$z������Y�S	��GO��#��?X��"�TS���/��:�,
�Wo�`h���wݷ�A�TK!�!x_&?t%���l_�����}�K��i�;|��\��b�v�O�]s �LYz�QSEc�m�gMw)���g�	�2@BUgQz��ư��'��o>'G<���.W?n���_*9�I�O�]fiE��x�dPڽB�նU��ੋ������j�NB�/5�yT\V��M�,U��E�z��w��6��z��v��3x^�)];_�k?��=ÇỲ���d'�`d�S�-�����ʟ�ƣ2��,ψ�}���5wR��U>[�ȁn���nN��@3�-�'�gI���B�>��)��D�LK�CQ�~S=z{W;�0:�Q"	��׏�ξ�KM��>�k~EG�{��0��d��7��Y�;�i����e��f]��s)(̪/ �Q�`GlYO�	�n�����!�J�(H����YOO]>�僜��`��Jx��@-gVc�����(=��p})窅��.�2B�SV������#}�qo-~�Ė�.�[�#�����a�l�*��W� �νXȾ=�[Hf��Z����Ƴ	YHgP:���?�:Drv �쬡���׼��^^v�EP+
�"�9L����Y��]U�g��!ȣ�Nc�mg��_�8m"�<�h4����;l����)a8�C�:y�
��F�ЈVj�F3���D�.YT�ZPԹ=m	��屆X8��^�f��&w!��@���*��8xU ՠV$A/�[g�׈Q��k�1������$��'5���)d�	{.�N��Zt�Bp@����v�LP�D����,Ql���\���qa(�cM�cχ��r�-C� aM����,�/m?������ys��S�Nc�b0��2���Yfs��_�U�}E9Pl�K���Vf�S(������'4��^@Sǋ�i�x�h�2D�|.i�$n�\�W�ב�ڢ�T��#�q.U��CH3�:i��J9���t`I�q��D��tbX*�+x56f�A��@�݀Ly&�>��N�򼴛]y���1ɡ��� �Ӟ�Ⱦڒ�͸,w�}L�rZJPE!A���E��m��5�DثX�g��"���%eU<��n���wp����Z�,h���p2��_��F3�[��mtq�S&|)�A����r����s�����j�f��+1��l��%%E�sc��o�Rz_ݠ�e��װ2&�a��~�R�M5��=Z��F�VS7�8M�}��.������s�h?�%�q������Lh@ixڹ����D�|!D��IK{O�5�]3nݞ�� r\h%� �.�c�@������N"��g ��m,,�`��%����1ɈN�T�z���С�ćWI�`Q��''�FLz��1 �A�S��jjb�Ջ��[b�q�;T݂#���uS��$X=ח�����}+��ꄩ^mV��������qp�/.,R�����YQ�����[	�ӯ��W�ϬO]ISߛbvBS���/i���(��ËEݥp��*�3� a|p�Rg;m�5���uy�PM1��uk#���ؼ����&{�d-v��C\�w/������'T�;�g-��;]�#���fP�<�%ы�ofW�ː,W �	t>��`�{�
��ptm�R�]T�����ל�2��䡩�4��������� ō�Fa�@�a��"��!wW�\B��u�`K���O(QX�%VƗ��U����Pyd� ���Fd�\������pO�@�k]^� ��RRZ�p�|��KM��}�`�bMQ�=s�u�JV�^)��s�	���Х���<��$��>�~�� $ne���4��lq�|����/Q�>~{n�P��i�1$\����Jvd�Wss4�m�6z;�;鈻���붯�Րb�;���6���W�!F�]�9�x�{��r�(��v�iu�bu�
�u��7}���P�1d�Z'�J���FL;^��5��ۂA_�O�7���.�$�lzG%ȣ����o
�p��V�wؙ���G��h�������	�}�
��j�>(^9�>�G	qG/��@IH�3~J1\��M:�ҹ#:8�#RJtL�H��v���ެ�I�d8Z9�\��� �b��B����C��p����Sx���$����G*1��ɼFz�ɅQ����&:K��6c����6	 1i�<P��k���K��\��C����ir�}�]l�Rю ���,��ה��{¦OX�cLKe2q{�M���ޡ���Fn�V��c*Jy���]�4��IK�8����L��=�4���6�nc?��R9�r�l��ST��#�Ѷ�b�Z�u�C7 #f�	�-��Ss��g�%zmad��t8Յο1���z!�V�\8T�"�d&���;)\!f���~X��T�>zs���oa��Ӓ���|�i�it3�VP��&�^� ����^E�3�J����W�'�j�\�iB�~��gb�t$����6)dG�1�c������ֶ�o��q��A�*t�����F�
]#1�s��Q�ɬ}�S̠�)�{Cu�d�ģ4c�t?&��v�!Ξ-���#������S���ΖR/q@'�=�]g`"�[?hgZ_���|�[�E��yHe�H����"�s���lÂE��+�&m��0>�����<�r�?��U�r�E��ɤ�"d��dK�8�/7cb��EV�8A��|Tj���t^_⳴�8��~˝C������nPF��mr_<v���V)2�欆��^?���c2;&�����4�o�Mt�nWA|^�Q�x��s��~�� VB�7���y�<m�oo�Q�ܧgvso�Y���ڄ�h��/�ۻ��eʑ���Wj�2���%��̱�K,�	���90�h�fR�`R<�h���g�_qe���.��3Xd�F���v��l�'M��k���$"4rYY��1��q��n*�	����Þpdo�W�Z �;��Bx��<��a)Z�l���"G����gD��`WU6�l���X��ؙ��<��w�V̨�j ��v�d�IV7&���uؐ.A����V���q��C4�\&QY筿���U��62НO2���T��W'�N�O�&[�/�}H��*�g�sZ�j�;L�۠L$��E�[���s�5��X+��ԫ;�X�49���R�6�q�TZ�F��#p���o���x����u_ǈ�ydH��ˎm���]��lQ-X�B������k>wL�2��(�w̄�Cr��e�9A��
���L�p��T�2����G�qHr�Q��V���2��m��J¯X�\#v���Tq:\Y���I(��DptO���:�B�B���47��P,p��7����Xm���Jn�c���+ʚ�Q"�;vk�ўW�H�{J"���6��U+��������곖*:<d$F}��^;�kz$iHM�J�R߻�Bv���L�4\�ۭ<��`lt�]�.vud/n=L�C����2|0-q`ma�~/��ߍx����/G��`����I�ʚ�����J�������I��V? �M���p[S]5f�B��F5L��j��9n�Я4�I�������i�>r4�D ��G5�ځ��W�v$}țe���4&���=u���3�y�[XF8;����>��~v_����PWP�).�h�Ç�;c�(%T R~�����]:�y�n��o��ﭹ�cs�t�H�w}���Yq��r���4�uH�8��~ʥ�􈜌���W�F�YW��Ë� ����=z�'f�N�|�̜*n�!�n���վTh��q�4A�=���W���k���Q�ٌ����HRrGP6�0�؊;3���ȍ��E+ y�+�W��4��B�Q�l�)�Un�@��f��ct�DX{�����o�� ������$������˂c��S'sҙH`�������� �\!�:�b�tK�??�8;�,��2
*GNg��1TI"O��ꨏf(b�� �G
�͏~ǳ�xP�oyd�ia�ћ��6M��pBJ��\O7C�W���|{�q==Mُ�W?�w�,&��OZ _���Tlв�f�i7߉��S����O!�Fl��d��Av*�y�K���?�@Gm���!=|"��gp�P����Nk��Af'���rN\��	��I��ߊ(�(�Fx
"�+���рj�{:����n�RTS᜽J�ñd	B�P�7!���#z{y�����Ćʝ���7�n���6�O�yۖ왮��9�h�~�d�t�ɾ߯�c�����7��g[к���Re�,T3P#!��t��ۦ>���O�]������'@�Z{7��1M���I�\�b��.Y8+D|P���.���1�9M�l�v+L�>l�-Fg��, ��q�������Ti0q���L��)����!�ԇ�@�� �y�܋꫖�Q
v�R1Њ�yˊ�HA��}����K����e�,����ƃв�.��n��bRl�G��h�+/��__�k�L�כёE�����^Ù?�Ɍ2;R۱�I 9k��G��F��F��7r�#���p�5���\Y�I���۳pye��H"�u@s��)�v��a����6����ÞA�&�p:����9_���c��rVV���D���!�q��R+�ceԃ?p� ��zl>j��m�!<ea/ ��*Ht�C�I-b[�h�)���qѩiT;�q�>]��d���<���(+@/�)�G|�bexێ�?S�F�r��C�{r`���KDm%�(��90��4tF�}<<>b}g�1���v�)�ĳ�Q���*������ ����Gl��.Ϸhn5<j�I\��p/�Ж/,A`�	���Ԩ~^��/�hpE���|9͹�S~��X�x��סL�>:6F�UP�hA����-IW��ί�쥍\#Xb�D�Kp�&�S�1��}lcp���Wr~`�s�+�����9"s-�3����S�#8+�-�|zūqz~�Ĉp	��Ϥ0�^�V������#����W�L�`�aA�j�׌Ɨ�1V>��I���{yp�\�����Zs��f�_���/��A���<�`�B�*�O> k������{/�G������*}ɠ��+���֎��.�n6���9�
}Q�����yK�r��&�$����ڂ��-Ӷ�ذ�EZ#W�M���Q:b�Y�D�������+��7]��C6)��e.�!`%獵��y��ꛕGa$cE�[iJJ�A��Z�>���7�t y���{��18��}5�'��W��!Xd�J���]��ͻG"���;�2:�Ǎ*3�lp���FM�6�`J�[mX�ݍ�Rۣ���9��K�z=\��?Uq�=�ἂAx�j�����	=�q��v�s��e�c�J�M�Di�6]�}���d�|T/G���9Č�̴	�����c��L'4>�z[�o��+6g׏=`�B̞ܕ'�Ҳӽ��J�� F�f=;v��^��e�y0�KJ��ð�S�w�Ykr9����lŹ�c�*Њ����Ht����-N��m�x���CFǖ��P��]�<'��p(����Dj�m
�R�hV�q�������q��&)7$E�y�� ��9���k�(�*m8F�TR	��2�͕n� �&�����4=��c�2���堌���qBT�`��%R�j���vQc>�'��e�JRPW�׃�A{�~J�sg^va�q�`~��2)�PUG�(��w�A"�.VБ�w���9��%�������!")�i;� �gy�b�.�x�GɆ�/���=7���?EU&B'/�e5�Ɔ|Tk�*�Ph���Q귓���fm�B���:dVIP4���q��j�᳐������k#�qjKm�1䐄����{��7,�6j�^ �
`��b��f)L�:�a�W��SG�pz�h��P�ق�>2���q��}w�:X��B�{b[�����@�
�0�ޟ��SK^�h�k�H*�>}Gu۠�H�<��5���s���$�{���P�A�ul6���k���P�p�dA����:fA*�Y��$�W^��>���	c]Ǿ}be��A�n��pb����q�*I��L7y@Ċ�b�ʂ�Vǳs���w�y�y�V����z8����g�0���4��@��Of�@Ϭ.ͭ}k�SCC��&�7��iC���D$�nL����2��^|� �X�y'���Ț�_w�eq���x�����He�5�O�I ��5�}�$������qZ�s�?��ɅF^Q��J�]qG��{��)��I�5S�;v�-�����ٸr���G�H�:^_i�������U �h�� h��nI�x
�d[�bx�{C 
�x�SI�℄Z�3���9 ����f����`��?i��9��뿃�5�/E�H�:��Ʊ�ԓ�x���~*1�i��Z�8�D��gS���F��zއ�B���K�"�#Ts|3��z���g���'%�fl��"$|�n��
�������Fi�#�>	DW�w�6��&`���3g� 1|#��߀j�b�ߔ�AzW�X��?I-&�6ƭ6�nPH�Z8S�R���E�A�w/d/�B�Q:��O���fC�íL&xQHl��OQp�S���_#3.�J�-
��������T���P_r�9��3��C��q�pC䣯����L���2�Eb�<���5�"���ڕf���2)}�{���N;�(=\�W�w1�	�2D�ʖ���$�"�p�A�zX���^�.�p��,���Z׃�r��|Hsӳ���C��W��9�$ҝ�:ܓfi�a��43��0 ���«�k�l4s� ��H�N$~sR����'K��@�1ϞH��[;�D������v�^��p�j橓7�H�({$�t�:�9����!6��qvUw%��+�󴓛?�8�A��:�<z�&�.���2�	>#u#��p,�ՎM�#MG	w�[���Ř�vϚEe;�K�8@�[��p�ＴHu`�B��՞n�+��JZGe���>b{ɪ�8���H𐢴�0��+|Ó�͹�s�?{�D{�1�؜�ED#�ʖ������m��]���zd�$������U�/.����"IA���Q/�*/o�6�F(�fbI�R��ߦ���$���Me�`f�6��1G�����dT Tm���ê���L��T�V^�Y��"�5�-͇/�6�.:�l�W��蠙L�����Ȑ��6|a ��5A�H��++ ĄP�(��~:\k��I��}uS�H���:��}�,k���u�Z�T6A�hO�*��͙���>��<�ƺ�(��S?A8��i(��瑐tU]y@v�#��)�1��th-�@�vz�{�[�m���H��Sh�˞v����oS�me�)�upc�&fm��yB��C#�8�s>M_�� 0c7� F�^$`��O<���޿.˴���b�
��bb�MeW�L��9�����E��5�@�z�gk�z	l@�羳��xW\��R�����T3�R���0i��*�d�׹]z�vB��]���H��k_S��FL��WRPu_�����lh�\:�x�3ԤLVu�����SqN�C��u�I�xAd�%�r�73u��1^��K(t���?!��`**�����a5(��Z����PԞ���	�6�/��!O���p��B^���i�D���
#���%�lff!�F�΃����A_�{�D�)��������{�8K��0s_����[��E�3����P<�t��yh�`�ry�'��	1NU����uw�}�D	Z�l��G�/J�:�������.xy��Ol���'u��'�⍀1
�����M�P0�(7;�����V-�[��d��'�TX��f�k�S�2	}ٺ_G�F����+[8�{F��6?+��D6�Ж0�f>B�ډi�ZpS�u��}�����6�� u�1��y�EF{
<���[-7������JĿD��,��g@����b�6�Ƽ��^�e��G$��|7��uaEfP�� U��濝�B� M�ɳ
i
C!�Φ�e�2�@l��AHߨ����*�3%�a�M抄��`B5�.˯����k�(��ׯ���e�v�̞i�V��������^W�vd�e��m_��j�}�p�,���;�7V]����^.��A�/�X�f?��	W��'Cl	1:~��/b��M���@n���ןϩ��n�a���S.��9�Y���J��rP$�6��
��2�'Cm�6$4zї��$��뀁�=R�\{������]���& W��[�U��;��a ޹��߷�<����!����Z �k����7�hkN��Y��^!l�&���Һ�� ��kd� �H��ƗNt6V�B�B�r�@%L�v��fPȠ�<��t7�Q�oZ��=�M��u�ttqWH���7-�5-����K�I��M��#q�ğs��3΋
�A�өO�>��mw5\�>EG��iO3���ׁ��¦����Y�<eSe*G�"�T��u��U��=�A(�6I���?�wL��RP����X<�S�M�����+�H+�|ٗ����\J��V�Z
O��a!�K00�:��F,�i�N��uHT�l6�zt �����G��4������b��C�Wb�w��ұ�����H�6����	QPdG�m��0��M�+�`���q�oD�։�M�����cl��Y�KM��D�a`B��
o�獦��{>�v���
�l-�ÞE� �\)if��%�q�RxL:�U5��b�n�������nX��M�CgĎ�������	��9��c����:'Tm)@����v%�R����Dd �`�OA!��E�RD�Φ�'2�5�`��E�����B؍�<G	��e���A:�D)E���;bPq�XO
�>�e6
a�6�}|�Fd�"���U���Xt���O��AT�u@ X��Bq��|%1�Fc��˷�vT`d�
�J_���+��PXK��3Ŕ)���`���<۩�o��7gx���A�:������M� �F���p����cfz�4vXw�>#ox�e�Wa^��i���M�4 !�����8 �9i�~ә.����_WK$%/$��ř�7�||m�ϡ�N��b�K�8�1��$x�mD��� ά���Z޺CxW�Ye�� V�E*sf:ԸD�Fi(�����=�BH���݇)���f��].(�J!ܞގK��\
�V���&���F��RLį�K{�P��d�!h�Ո������0(�j Dr\M]���	�?�|Mp�y��xD�Fg�
ou��O&&�m��]�����������%lOӭ�ogh�9w�]�䁤����z�5{l�꿝�j��c/�Q0X/�l��y� �l�ŀ� e3D-7�6Oy	:�-� ��uA����.�~p���=
٤;%JA�dW�Aƶ�Y���_�c@��&�� D�i�w1���-:;V�F�ٰ����zs9JB�-���s 7
���x,?�$�jO����0;*��qr����y���D������=E�BS�bUb̾*�Pv��Ր
Ya������E0F6C
�R�F���������+}�V�n3���M�}����7�Ȟ�x��Xsgz�@���d8�t;���	X��
��8��<})N�͵�X�Ψ9�f���O�wh�1L��8�H��Fޛ�f��%&J_[��?�o��	x&,i�"W^���a#V�РM�6X)����ަ��?K�T�S��R� BKв�o�.J!r�
���5ܬ����	�u�lh���c���l:���xQ��"��P?�씆s;�O��Sf�F��n�mQ�F���\@F�LI8�b ʍ*�uSC���~ʢ>��ʃD~lsO�ױ0W㎭���nQ�p�n��A�})��YE���+�1C��-ΘA"mX%�g�o�*Sq(#З�~}z�Lˑ���,�43�c��S����,G��_�+~�+��9�J��k|h�����������:O�K�}W�<���/��Z?.�eS���ɇ����+I>0F�Mc���nUB��K��*;���R�Du��9�J��Wͬ�g}J���2�G�7�L���4�x�;̶'Q@L��R�J?�E(RX��"���(��tܜ:򖙴�rG)�4=��Ķ�₹l3���8x���PrxE�/�$���8�11U�� ﾚ:I�ȶK:���/�b���K�m�Jf�-�y��0�Uߥ�9���91�.Ԩ �<�1�rU�$B>�:��֟X�k��C����;m�%P,L�32�-f:>ʈvwO���Q8E0?:iEfQ��1ҧ<��]#H�!�@7��1��1S߼�bU��D���{C�B�_�@��`|�C5:1�6�͔{P�#�tsz5�%k�9/�4˳Y���,�/U0�!�UF�|�$���G�&��<�7P��;eeO�ʟ��f\/<tX��?��H�2a�,?e���\���������a�����B��٬�~t��/���=J	j���-��g?Atw��������u�˛V�\	�g�GNuE9~Fq�pW̈́Θx��J�QY0	�� fn�NN�L�0��Hk�1������GokF�{��;�Ư	z�?���E� ��\��-j���d�u:3�[�9�qL&j�1؁�N�d9"���:#oq������ezj�X��[I��L�jn�8�%Q�E6Dc�qF�����a[��T�6�Ur%D7�<��t�8l�6LP�_�;�]i��B�g��f�*�.��(�m*��,�<����W+�v���*�¸�����p*���U����gPdv�k��.l�GݨC���x?K�IM^��}��������_WW�4�'�v�:�@P���ɢׅ�Z�Ɲ��&�)�+<e΁��3H���ʎ�8�?,�,�hmkN��e��� ��,_��sTdi�Sc=zz<[8����E2����=�+��M�-� �2��~b��������~�������-�u����ڶ��}Z~Iڋ�vK��K�P�������O���B�n���ե�s�jg~T!U`Q�EJ�V�_Ū�Y�4:�7�8?�%
԰�	j��qAOjB���� >!&	T�6TӦ��v��߿�

�2����;p �VLu���U^T�˵}�T���dˮ.W՗�t������0��u)�:"9Z��Z҉#�U���
5���X�����F�6���0-;`$�B1x>3N�d��{�r,@i�s���!K�J�O����`����#��"�wf`�Q�N�I�&9Pn���%��Q�bxd�ץ��GWwf.W�ƥ�cq�`���@�<"�"���}c>�I���/ML��L�Ԝu.$2H�Q��N\�'i���
iV^V&�`�L��,`4�4X�a��O�|Xd.�!�����,��z�!��]ソ�Bc��we�ʥ>�Z��#��	4}dɐSyJ�4���!+�?~�^v�z����ϳSי�V��C�k!`��m�Q�� /����X��s�XO�GW�v�>=hHԮj8�Ή������i؅*�g��A�[�.0�k�p*��=��~ad�U���qu��IhF+vh%���,��8e���Y���\1�"���5��R���d��R�����o%1�o��l�L�*����I?�}N/+�r��۳�A�?4gOŋ�\糿�k��)d3q���(����^f�[��C�B�=�ح�G~���v$j&#��rJvM�N�r�&�h@9n� W�;v��P���^p ;��,��=���8P���tG��J�
'�`�y,&"Gu2Lf��fx�λ?��˂1���>���,�̏H�#��1���|(�	"!��ld�'���ݐR�D��=\�NQ���}��wG�����R8H(*Uq�\����w�9k��ɦ��CD��nq!����	a��)���Ȗ1?���u&��?�E����qio������ä)Q��0ԍ�!X!/(ف�Ga��D�@A\�ر�;N��Zx<%�Gq�8,�M�;����6=�(�aX�yy|9��d��U⸲�u��3��EھHI���5�����t�빶�ь�'I���9��m��s5�p?�z�]���{��N���3��]����p7�l�4e``1V���ȏ�,\;�,���J_�����ovtJ����Ӎ��D �E16�6n���zUys;H��r��n�v!ŧ�醚�7&�Z�Ev��]0"}���#/$�BE��ר@�Wn6ڄ��4?�Z��#/  (�8J/�P�_$�yZ���nY�"�T�7��&P�����P�jz3H �����	�+갓q����)�*�7��$��3�h^p/D�Ӵ�-'�f3M<��Q>����+���ՐvG!P6�)�mq�����]H#�ο&��߃��c���b0�V}�.��m���C@_9p��x�{�z�T>/dQ����Ll��\�LeL����'��#��	uD�Qz��f��b\�\X�,���ӓ:?��Y�����+�Q�f���q�v�	�RG5*W��9�8���:��Z�����)�G�N��:SY��چu���@ESj�)`��&a�XX1�Y��؟aY����nY����#P�{�\(>�g�N�ƿ��V�ݧ����=���_IR��a�+3�a&�φ������H�`�d$�fs��/��Qu���Q�Q����u�_HH��NY���߅�6���dyG�z�ԩ�;#I��j�������+ wA/J��o��GM��<���L����R��m��v����y/�l�X,�L��� tl�#��ɖ���Η�v���ʕƄM}�o�2��s�eL�y�L��fIɣ@56��-��Cm<&�jsuqq�����I������wK�e�V�KE��ڽ5�N����
b�����G�X�W���L��k�Q���uo^��6f[�[�)&aB0������e� �>)/�Gi�����LƔ?W�j��CgS��ѷ֐�)a�.�xn����!	Z!r1�+���������ɝG�����:��o32�Soq���` �A��7s�X3��P4�1�i�m�~o4��&J�����l9Bi�[B^�B�ti4G�@j�p�c|!�o�
���P��iy�=��:�t%z�Ş�Z����#$A�u��1�<BL1a6ֻg$\5ѥ��3��=�a/5F*4�99���kl�B���E�C!��e Z[�d�\�H����u�(�Ԛ�B{�tȡ((�%M���i�}Dhuᑜ���\hSb�.��V�V��A����O.�`�L7�qOl�RI&P6_��k��hLgZ�n����L%9uYM��?/,���WUH��
�b��4��*����7��j�0xRL�SOHx$�ާ[<]���Q�5��� '�?��JOs�{$(��f+bgaj&��Kr;��ёdB?���	�y�u?�Dܵ<Щu�I�n���~K��r_�G;X����3~��yFַ�(�{���R��A� e�Scr1~�W*�L�"w"n�hw�,J ƸիL�b@�j~a������kB}����PQ�!:f�؆Ш!o{�7#�c}e�מ�({���d2���j�I�O@[1|6U���]�Ͼ[�A�s�_��xc=Փ��		8��c:��c޳z}���nm��1`
�:����
&�H
7�����3�3n�~`T�t�3����ḱ�JP)7���L�a�v��t��2�������Hz��mw�&�B���ˈ��j֚}Z>f�Z� pZ.K�vQ+�s�����o�#ӋANgf�DQX ���6P3�s�қJ��<r�2���$�g_����x��͋�&x�m�|ʳ������.1�&p�g%�1��4����0��tu�	�ָx�i�����Ќ�V��*S�>.1�ƥ��VA���$�?���I������s�`TYJ�o����C[:��yk�T���&;���Ӎ*��l�!{(��A-�:0�3_@��# Q�1��썩aA���0���lH�_o�"�ak���j�m2Ҧ�P�,F�$�q�@L*�r�|C�����⇆
q��<C���z2�KBSK�䃣��AX�YnChN[�fȵ�e�7��ؗ�ӣu\�'�t��&�Č�,�jҎY\o	�N�.E���m95��"q������J*�qr�L�]�gr��:�)Q�z�ٙe��\ܠp�\A�z\�	aa}����X�Ѯ��� ���n�ZJ�=җ�TB����1�V��Y"EsP��2=���V����,Ы�kG�N��9�꾸�E�4�	��x����i��D�ܓ���R#��
z��In]�>���\)��\�u4G.M9Fо��L<�lO>Eܸl�F���g�h�I��X��ϻ�~���Wl��%�[EF�.�h-���;n]q�rY8Z4��2�@(QPa`�������#s	b��꒻��(b�}W�Y�6�d(;�P,.��h�W��+��$>�a���u��J�d�V����j�� G�[9f�򽟊�8C'��	e�ę�F*f�2~K'��_�D,u^�C����Id�-�$�iQ*1�3GE#u��w!�'��\���~�~8Ŷ�o��M�l�1Y׌j��W;"9l�<�a��3S�Rz�_�ճ�*�[���Lq;�JZudh��/����z�@6��T�ϟ���\ �/���� Á�v������-�(�w5�M��]a�	�0�Z�����n�Hy�fԋ{�e
�@M�q���f�6�@�R��޾"&4�ǐ'�>��r��:x�5ڵN���<��� �Q�>)~hv��2��^-����`(����ʐ�Eϵa�,��w��Y�_�	�2�mH@�雮f&/��	n[C��`dO�执]���4�x1�<�/L�ӣ
.���(��Au�۷,J �R�R��xϦ������q��������=��y���5E0���� ��ݿ�z��!�`[<���쯂K�
;�6�'���6���Z,�v�\}&��:ܷq��;�#=��I2�<��`ir�~�.� �)mp���Λ��O��-��O� ���;FM3ns�/���\��}�ַT-�I�ԊXж��|̓C
p�m?��2`�d^�������/gQUb�XC��i@0�x�b��+�q�^��0�qx���Xˀ��IO ^�D8�Y�w-Y@cZ�����T�B>zv�L�?�-��Ƥc1:�=�pd���#���L�A�[ +�5tr�qO��4>!~��
�֫�F���҄�J��؛9R��M�������u�-�RD��O�a��~�`n����ۭ?ϱ֕���K��Y�T&q�բI<6�wj3Ӟ��V�ە���"����XJ��c���c8WdՑTv��U�Bnk��p��:+��M#����h-��za�=@�o"�0��vQ�M8�i.D�,������	�{$��G�R-8�-	�B�K�SD�� ђ#�\~_W��,�0`�Kt�R���b�d��6�t�'!�A����"N'���T��I�^���%O�hR���,8�Q��,[ތ
=��Y�������U��Yϵҧ6R�u{�4Z6��z���qO�
��a�;��D?{)IX�t�c?��䘶���g���O�x���4�<��=���ro�m�m��7�H�7�͗gq|�C�w:�P�'��Onq�k'bi&%9�O%u��mU749-妽ǹ���}�YcN	���'�L��-�g�)����������L=����Z�<Ю�S�fOa#�<��1A�n��`p���e�:j���tYYz-��������)Y+~�!�0�Z)��$>
��i@
7�Gɱ�a%f�'�Z�ňO����(5l�`8�� 
����z�.��[5��HI�l�^pg�t$��7#z(=���r��s#�15&&aVն��3���sG<�8u�L���^c�a���"�����IO�}¤��R�>�ވl���|X�z���Ճ�g6�TS ��8
P�_U��b���ʟ���]�(2��o��D�Ѿ��.,�Ơ�Xq�~Z�qh���5&��k͞Lk��e½z�T�����TK�!��h�9��Q$��<�s���s=������fӿ���[	��fT$�tb���M�8 oշ�耦Ѭ�Wj����/��z�&f1IK]DT2�7�Ѡ��'c'�O4��Z�U�HP�5�pp���`^��I�˖j�����j\o��D����>U6z 5c����O��8#Gd�hPuy��x�IQNa�)��\Z��x��Y��"}Y�| �igյ��i뎽 ^7�	5���'�&�	�{��4�b�9Dws���Ƀ)��n�6��cɡ@}��|�	in��R?�2<�����?Feu��X%�qo��%��i1e@�Fu�K̝㵷B���P�E��M��h�.�=Ѣΐ�$.��f�֋a�3d��X���@�=�_���~�6	�n�ܲxyc��	�����$�I��@U)��躂���f�{�}�5ǯ֤�up_�jLĂ���S˙�Nd	� F���dn�M�A�L�̱�с*
\B3�/wIVy���J$��d}�!F�����w �f�4��MD�|@h�vt�ʒi�9��D�LU!�f_��=w�=�O^�L+������b���_�� �C�B����@��G���.�O�^s"�WN��q��A��ϓ:\'؈5��%��{N�Aq�Yc�^�0�p�@��b!�g�ՊOn
�2ԁA]���y�/8�X�r$��f�g��_{��A�E^����\1E��g�nb��@�ʸa��  �.��-eB�܏TɌ�&��Ԛ�Zoy�!��0���k�4��\�	��K#*�-���c�6��ݎ�U�~/��{|��Nk
F�'t@�a:c�d��W�NzO�sC�Vf���Aϭ��� ld��U�U�����t>�7ܹW�w�$J>��F�O;��U�z��I�y�T�DN��tg^N<*�sٽ��9	�u��ŕĘ��^��&�6�1��J���IKBC ��/��\YE�֓k���
�f0 �u&���6� ����6+A�}�e�=�UR�.�@�&<e��=lR4�w��+��U�Oܘ����K>	r�m���ˁ�F�b��P��P����E9j��8����!Hy6��gs��B��o��s܂?�J�=��Me'I�b��`iv�j�}�{4�E��Zmc�{����2"�~������xڷg1uǥ��|�Dx}��A�_szܥ�I4Dzh�q7��6C�$��� ��P<��i !υ�����b/~��aX�(r��j�����B逄C���
�ת��������j�DJ4E�c�����$Oc�ܬu\DO>���T��0����v-�]�{�K5;�R��LM*%�l�Z�I�)D��:��r�I�Ӓ�F)v	�T��Z���v��X;3�G�<)�=����ړ��/�`� ;�b�m�P�d��#�dCS�����V-eu�4U�dBʧL�s�(h��[�Y!�8�̏Ɍ��G]�g�[��`��e�ۖPܑ�A��!�}]2�K�4}X�<�:>/��~ͬ��nY[_�,)-B������H*�>Ȁ&��}#�bwV����7�1�XA�qh�,��c�+�u�_I�t)p�����*(���V�U�gS��/ʸo:��h�T��?ag�Lё#&h<'5�&�.�=�����X��&��jZP�}��{\�?��&�ԓ��A���;�������J��c�����đ���Y���`��^�x�2Hry>�[�<����I&�=�W�]o�U�<u�n�;�T��Q���[g���t�����IwC�,�]����*���t�l�-Y����B�F$��v:4�M����h��НZL��Ba?���ye����������@�>Xh���9r<�A
��xb��$������I��̏�"h��2uEp��O2�6��i�|y��=��=������3}�}2#���ɂ���&[�=�5c�
�:5�ɞ�7��o��76���/����oz{�c���t�ݗ<���F�n;�C*#��h�i�r��,/�~�f��Ъ�e�\
��	ʝ�k�g {�v�:��9}��+i@���L8s�l�)��&nni<�?@��bP.ڥ�_���J�f>,�J�B~��!D���%�Mh!�4&O-�s���_����KFQ���z��~�xl�/�y��E�����U���Č���X�6��W�
MT<��X0%cZ6:;e��g��YܞP����Ag��T��:I�g�xYђ9W�eR�ᗐw���0I�$��r��n>y�G�<�g8RjPB�>}�HT�C��9����f��ļ�T|H�n%�ڭ��؂nƷ%a9�6��N%=��ѓ}4� ?!	F�(�ZZw����/W��;A`e�7я`��Wk^]����PɻFV՟.b�[�����M�GM�u��UG	7�g�.�Һ��I+lɞ3��crg��A惯EB����rFz��4:���Q��-m)�]�?�����l�]?�D�a禓����dG�0�;[����I,�=�k���2�X�F��ث��8�Eb>l�H\�c�R)�*Janl(�SpNUEp�?w�H�c	0�y�k���i���]"�5�n'K�	���K��Cݷ.�s��Y�!�;�ߎ)�5�+�XTOy�S��}�QС6iu�gr��:y�2(<..DPv�d��t�G��ę}�~��4��Am����m.�u�K
Nt�.���p����K�z��N?ؿ:C�_���1\�v� k=��8�iЫ�Kx�	�
��0�z�~d!��l��`�%q��ylI��>�GrԎv���tt���ҁc��hq�Pnh}e?FC�?
�B�(�Y�T֚�'�����3�׫��p�z0*s�S9�S��.�9W.�5�l=a��Q �a��Y���!�e��.}��Oz&�"jCPT#���.�Ǥu���/����<i�t���������t :����M�P����
.>��}�]i�fC ,�,��M4;�Nq�=�MI���e8@�Y��z���.�Hh�/����_��s��M�Ïy����5�hS�Hj+����K�1DwB��yD;<k
�H�ݘ)g�z��;��6�i�}<�i���j�`)�x�?O�u���^���0����g��uUjk��I3�!c�Wt&fk�w#�ˤ���[q��M�����u7�J�(c�2�	-0���@D0
r���I���d��iC��ވf�2y�t1�Y�d�}��`;3�^M����`p= uã�4=��r̫n�$M�YR�BqM��Ζ�«�٦��G>K�:©U�?�J��d����q�HO��fK0\��ʛw�2��7=�w�D��,�oT�3^�.�T���*�&���C9]��'��s�T=��R��支���`��8=��/s@:x1������f��1`;��$c�;����m�w��|�Ļ0�����U�����<��9�3����ء���oU��Ʒ����*�
����z 6N�1��qR�����eZ�gj����ٶ1�(.(f���^�	5v�'���۬�P��|[	
�{�"m�HFE�C6��3֐ͺ��(Ԋ�X;�4�	3D��H��J���/i�2M�ik@_�#��'����. ��@�B�`��p�zC#�n�9��A��Z
�L���hbK*��r�ɅYK��	���P헌�p	�
�5�q���d�11q�;6{��� b�C���n�>���g�K�k�+hu���~H�6,ԕ6kk!�����4ZYn^�;�~dݰu�6�J)�-�T��6ұU�OE7�_&T/���`�f���� ��4p���2�� ۱�ɍm��"6�����e:��8�9ވOz����eq4�0�"���_����"�)�������澔٫�^4�u镇�3! ��4��U��Y .���+sAI���4�Q)O\o�V��|� �8���s��k^IKhS�RSJ������q|}��9�|2�9�K{W��	�{mw�o�Ť�E�.oIM�%���R�}PΎ�$l����@W�����ϱ@n|vQ����������'�4�� �D0�5|��d�1֭u���)}卍�WǬ(��O>�'�v��	���ߋִ!$;�V��;c�@�.����J��+�33�*|P��)q.�tg���#�5�Qa�%�Gt�{|���J�FͰ&Cs��O�5�o~�AϚ h�r��I����X�i���@h^�L[�U3�=��� ��M�6��#�����&�1i�j�K�2Gd5��	p���x��l`�������D	��46���֊{�d�n��bE�����������CZ��z��N�E��d�ծ�n�S@֜����~)�v�{����*h~Ŧ��9���(�+"k��sBa�o��H�����N���oUXLn�kO��#�^�"�~��`����Jkkq�˒�p�$
���:-�B���0�s�8��3[���b�Ӧ�����1G�(oI �P��A���b��@z��isRl7S�� m�;��4\sH����jO��Q��j���3yR��1K��}����^ ���q3�����@ϗT�wfo�����=�h0�_�[A[�M���gu�7�Cr qA\��O���8�)|X��asT��{B����3.(�i�/��EI-�.�լsE�/��22���Mr-KY��D�.��^ZR��w�i�q� ���/��(L+c��
L�L�u쉩���>��q���p�~��Ԁ����e%���&��垙%��b�¨Gu�.�xy�x���v�|��\�{��"�����*�5��:����g0�0e��� |T0鸲�m2�e{ul0g�E�Wta6��Hbq�|�7��/"�G��+��)"�,�'���cQ#ի��G��������1�����c�6_� .È���&����|����"���J�uv�E�
�e�j�4�u����5M�R�+A���62�?���"7No����O��3�ks�?�Z���_p�}U�L3&5-��K�w�2�T���a�NL�R�v5l1�[��X�t�q	�_�_��~$��VE�i��P�g#i��x[ԝ��|п��N�4�B*�HD�6T ��]�5�0ɲ���@�l�إ#݁���1`8#�Yz���\j.��ɺ�o�,f���4^���}���wyh+"n�,tt�g�#{I��?���8S>��/te���;�9?4D��K�(K��<�g�I��_ӥ0��R��F+��*5_�H����aw8Y��vqP�9Vs�HU����d#ۖ��U�%n�R��%e�\���� �.���qmp2֗<`�V��{#�ȇ"����6Zk��P�Y�Ɓ�P��d,{��矑�)o�?�� ���o���WX���y���C�����M���T5h�8���:��-�O���Z����:��Չ>��m("*	��v)�^_�8�%~��W��6��[A�.���� >����5?�G����뚲�H�o���%W����UFY�j?�#�q�"=�p�_�Φr������b������vU�L�����^XD���ξ�܅�Kb��h�[�ɋ���~v
H��XH�h���5�C˨{b����>?]`�VK�`/�E��N�����lӡ*�W�Ю�Lݝ�"�QB(����3.��;ޛnt��Cw����b�|0�H�*>�5����d�x\�8S)~}��I*+͜��ns I��wq��4�g#k���f�~f5�.��i%b��W�ُ�;Zy���^�ǣ�����Fxh���A8�0��(��� dc���)�Ԡ�ʔ*�	�w���4Ow�1b�|��yM���� لY�k�v1jV8�(��cw:�y۩X��{,#�1w�$ؒ��c
���ύ��p�B���i��y�y��>�. n'��C��ĉ0���l��c��"��X�]a�i �\��z�pj�f)\�S���o_�w]�r��C(Ӭ���#ɤ��@��!!XE��e���|�N blR���Z�9pi�5��E\-��B^���nQI���-2U��:u�T�Q�S���Ϥ)B!\����7v�'�CM�C%m,�'`�W���'uBO��3Ρ�[����֎�����v����7�7w~�1�h3q ?����{LI�Y�.J���ge�(���a����0�d
�#�� �nB�M��nœ�&�K�k���K�p�R�tA��������kԎ�Doz ������6�J4���n	SF��W�jЋ�k}R�@6�R�C�]�� h1$9`!0	�`��栜�J����)��:����?�a�_�&�d(a��[�eCUJ�b�,�	Ե�^S!2�@���-�%C��`����4�pU�_#_E���L�.x�'���q'�j��ST���{)�I���"��? ����`e��D���=Vh%6	w���߷[7�1�c/}�q����m�sqP�4��Vo0�<`V{�}�֯���5�6Qʹ�/�5�g87yĹCH0R�%�ܐg�ȆqD��\�)�r�+ǳm:��� @��0�f]P:J�>�$�����]��y�(!zD�AJ������3wp�m�jJ��������X��} ��&�F��	�"�}�O[y�(�@����'v�wP��� [j��	��k�U����K8��]�x�޻g^�����j ���exQS��C���b���] �f���d��p��A�a�<����?qF>'5�:HS|�+�w�g93��k��OJ�X��3��&���W�#X��Jw���	�p�]?A?��^��@N�� P)9.�c�F n`�v)Cn���V�M �1�����5r �΄�/���F�qFg�j�]f�k�-�e~'�9S��,_Z3f�{�����E_/�������Qg>���j*_H��ߊ��>�"�2�R2'fm\_ʅY7��<;x{��Q*�nĴ�nqL8�&y,����׋`��Lkd���r�D���Zz`6
���'0�:�~Ha\��&�CR���N��A��:��)�$I�`�I/��D#�k�4!/>[K^�S[�X�6����vz���Cʇ]n�5����MO:����C���2�
�G�ZX
�kYfp��Z9i�A��M��>߽�r��7�����۝#��~D؁=Ҁ�L�d?2�ߧ?8���x��}�{%4#�n���bıf�Ko���{��×~6/�X�O�R���ߡ�1�J�Cc�'��>�O�0�9F�}RFo����Ӛ�+:]<+�=��J�[��c{+=�$ �?�FL]�<�T[u���P���ɡ�E0���	&lxeB�#���ب�U�D�-w�^�c�vc�������Ilk�)�k�ƏQA���5�c��/<�
��Ko��6N׆�]�q���U��tst����4�pI�bM��3��e�LY{ ��Q}���B=o�v �Ε�<���=I]�[c�{����Z8����'��N!�
dl�VH[�ߔ���MUH�_E��	�����Sˡ.}yA/�.D]7��B�3eN�����GY6ΫpW��PF�R=��rS��_g�U���C���Byp	ݦ4<���B�3��D/�Eo-@��-Z�6+rh��\gc<�3��B�խ��U�W0z����&�����{���vu.,ɇ��pX!-ܴ�'ܭ�.�
H�_ $݊��p¥�	��;x�bCfH#�	dt���6Uo�������L2*��]З������0�Gi�
�`}�8�#w�u%�~�7�9tN�g����~�d4ӷ ����4s		4|��N�}�'�Z�X����\ĥT�7uӾ��v/)XTߡt��[r桭�6(��ф;���-ߎ��9�_�2$��v"3>cܜ�r��(�,I��>}���ubT��X!��V�
�	��Gw5M��PDJ"V̜��E�@y���6��{��.��s ��b'[V��7ZV��0��aO��?��*n���Kؗ���	��",�&6��l��˨���E�IQ5�쬨�+*+����	�q��?�mR�S7�yZ̝+F�f���]?z�4�L9�m���0�o��BLqSC_!��9����0ך�d_UX8K�;�k�~�7�Fn�@1
�g1�a������TE&����1�&*�{���g�=�fm���szYϳ��ߛ�"�h�"H3�L"S��23���P�g��Y��o�O�I]�O�T-��@�1ŗ��=�M��N��x���h[v����,n0��R�#� X�tލ�=Vf,��$C:�f�g�c��fЎɘ�j	��J�<hND.���$jO%H�Tǿ����q�f]G�]��9�+������>���m�g;�Q�ifaK�Q�h���}�dX3Y��6���@�s��f�p��L��{F�����SgK4�������k݆#�8>sI ��c�iG;�H<]s���G�h'Ѧ9|-8>��5�vh�u	+ X��>eL��
5�I�����Ų�JR�e�=cK��[⸴���e0�2СV1���	Ƿ����2`:��8I5������:�1zOjG3S1�p�h��nT2;� ���2�cp���u���D�K�f���`I����!��}bL:4���^�IҔ1��W�&��(��]�����p	G��+�kd��`Gkz���f`��+]�\�b�pp��'f�>
u~�H�=+	A���B@&CDa�2��gƈ
���`���D����@�8��,�8G��^�=�Zkc��ņ����$ ���*��{|����?)q��a�qtɕ�0n1��U��C����3�n>���8D	���]Uv���>��lL��g"ݦ\���8>ļ����h��t�Yq��"��b�'���6`�?}L���VOߺ�w1{�@�b�0��w�g�)�×q��v2�?�]�a�n�X���G�gظ'���$��K����������/3Z_��	����;�b[(�L���M �"���3$��B����fṄ���X���oD�V� �#�1�g��_���	Q:�,�P��$)[X��%3��,n�	5��1߉LnU3	���2����S}��;��ǐd�N�`;H�������~��g�K�N�.����g;�H� !���iuzoD�����O<�����Pe���QG���E�������H�q��mIQ���%	�V揄�����;��S��l�Rp���҂�(n�#|oe�Q�	b���{Ӓ	��hN��H��q�&d�Yt��>b1٠\�Z�9�{�eV��d� �t�WU)�����Hƅ�g��C�����P��=d�*2��d��?'o�Ѣ�*u񉙯X�ʺ��Os\
��U3����9$�m9͡)5��,�jQ�Z�q�2��M���Pڒ*FB_6��,I��F>�;��ϕ�������	�b��
.�I�
qL��Pِo����&=Y#ϕSaAgg�WǴ�X�!�����H���ð���A��x��̊�U�����C2]N�.(נ<z�F��ҏ��9fWgE-P��||����RLeH��OA��`�j��G�ڣn	�v;썾�r�x�Ox��g���[�+T%v�B�A�33�?ʼn�\�i�����>3f�/�vP��Ɂ��qP��M�ʆ��*`ob�1�&V���st)b�]�ő���L���fՖ�'�F1~Uݺ�\�V�̓r�����LZz��t�x�����A���7�E.�h�5~�}��]%�h�m�i!�,N�p���#Q^w��:����N�t��][��q���Y�_���}��CI�X�5:u�K�U/a��)�>�¾�~Ħ6�!������ )'�Ȥ������t#�UH_;	��L�<v̼�(rd&�v�Lr�O�v�rY,�啍�F3"B�=�T�m:-��ڃ���}���3��>��X�y�{�d�>��ş���)���+ž*{�EC�P����	�Be
�q����O� �B��N�09Lc��jЍ}'�|%�h��2d�c��&?�o�p�#f�`]�3nC1��n+O]F�>�:m�e�)h#:��>���1�%�~J��������b�;c�,�F��8g���܃�`�;�Ůb  L�*|A�@|�>���C�ak�{)\Q���g-6�vk^��մp��GD�TA���F�K�á�)m�x��'x��!m�X��x�°��0��9���<�&<ܺN���	��J؜�-�P2PJr}��9�D��t=�ܻs��,�'{�>��{ě�*�hQ�L=b�ȟ/������'��y����	��j��³0BQK�Ȯ�"�Qx*�d7(����B	|4�f�3���^}-W���⥽{q;mzL�d(�Uv�.�S��Rz���aS�36nEWq8��4�خ,��̖S?��_�o�;�3I�9�3Eˠ��ٌ�VL�[r�}}��1�q&%�cWb��F�ڦ��R��	���{�hM�O�t��H�х�o�)Y���h@��܍ ���M#���g�ے
�`��瑲�����-i70��.��i�����"	e Ds���ؼN��y�#U�Z�?�}[�s0x���,}��Ljm�T��zi�b�:�.Y7y],�E�Ϲ��q�K�v�	|�$?�)�p5�7Do��D_��:��0d��K"��w�P������B ��ܑ,ndS	$75��bi��@�6����/?)�JĹ�!r i}|/zOt��=$�ʉ��<��Z�� ��B~r�9��&ݎyO�ewR�Ej-�/�����|�~E@�滢X^P���\X/py =e$�|��+�\7#���_��:k2��"�'{�z6��ݎ���U����[B��h��jE�>� �2��Wt��8��Af�S��5� �c+9�>2.��T�u��X��cl&��^�շuv�ϙ�<<W�_(�xC?Ȟ^�y����� em}���ܒ+�dg�"&̬�D4���(}� g��?T/*�o���Q���q�����/Ȼ6v����[����L�xܾ�?O��@�z�.K�έ��U��J�����"_&���t>Lm�qKK�O=e�D�ɼd��v�*ݱ^]XYWeJ�)\���*c= Cӻ�Z�aH����p菾����-^\�f�m�gQ�HF�m�H: �}Z�t5�����= L���F|�ݍ�7��y����m��~H���L.�ǻ�2���(x�Е%A�T4�7�E��Nh%��3Lǯ>��f{_#��n{�Aֿ��t�{L��>cE���,��$B���"����W�H�ǭ6Q������ʠ.���F�?�����ϧ���S~ *�������D�i�r��t�G��F'�Hf?�d���;)?���Vrii�ǣc�w�z!�|)�Pg����_�n��L��b�=��dk��@~�5���9��0v
�|��"��ٓۮ(FfV�-ʔ͖njp�e����ae�+۵P_���v��\� �.9P���҅�g�@_{�ɒ`���}O�&����*�e:�6���2���(r{
��Q�C,����B�ZD}�FDs���.����,ӣ�]�.����h�K����VY�3���'��Ug��㚊���"���El@��`��8���
 ��"aZm�4LwTW�zqB9ij{E��C����ꃊu܏�~�����}��n�!X�+AJ���R�	�ykp	;wnh �<����s�}Uq�����4�<�XWgVf�g����p���TR���1&(�h4�gF������kl^�����F�£(�6�r2眙��Ъ#�^>[Yy04]M��p�GB\�Q�>�G�����C�"��0�s����.��íw;�!�0�M�\�a��J�ړ��ɕ�>�>����ᛯ.�k&���G����^T/��(��{_h����)�|�I�Y�mvI�+����g� [\1K@�U)6&�!XD��ْ����Oe�-��aM���ܩr�!;��{[�L0���:�n!s}2It�j���I8�j��CO��yC��.��o��H��j8����[�T@�4S�n[q�\��Xa�(e���`Q�7@�gER3v4��8<R11��4�O�L��N�ѡԪ �7,Qy�"tp���&��F
��߹�.=�2�-ԍ������⌮���we��}<����E��}�G�焠h��K=��J@wۻd=��E��{0�|���w3�3�<'G0�Š�0+�K
���.��kj!RkVװ/��ނ��*ݳN�H*��IR?k�2�o��\h���k�I��;I��/��'g�Y��I$�	Ay e��f�)����0�$�'�!EF�c@��T����|��1�S �<�������lN�MfzɊ]��Ky(|æI/ږ�{t���{���@�^�2�y�L=�,�f�Ө��Jͥl�nGw�E�_cr_e,*"���[��lQ�y��������}�?�X�/5`� �I"L�t��S�=��Ҧ�A�g�9��Fl_�I(�KIh����{�FS!���o�]�߉��s�&�{j7���%�˩��Ss���2��h�AW�b��{yY�7�F��Wζ�cnE��2��O�x�5`2A4f��������� [e�%3�\�x�?���-�Ҷ��:��o`͢핆x,	�I��K��3�ؑ�(����T�"	k   UԤ���I���:��˷�\\ؓ$�Iǰ��������F0>kw���$�ҭ�z~\d�e�H��V͊zR�p��=ex���Ϝ�0��N�[�ؐ) ����V����?StgW/ܶ���)��,J���Ƚ9$�}a�;xF��t�����w��uO��؇�V|&��l�@����<��e*��.��}z��q�r�x�M���U�@�(��_�=�3l�"zE�����jX�����?ѝ1���F�`oX��õ8Rw���.a=~-1뚻�IP\���H$eJ%��}�D�z��G��ƣ���Kt�`pV$��GI��U�[�כ���=��<=�l�E�x������V,��f���75�J���������gE쬰����#(_�$�#U������b��?J�c$�wի�Рcv7�j
�Riѿ�K��O����E��=����2����u�}?h�g��l��>���ւxX֓�5u�=m;�P�?)�y/�|,Ǚ��d�[��U�kql�!��[������ �r�K. .���V|ۨ`e���DDc�.�!2f��Ҫ��Sdק��|��S�����"�Fw��~���{��J��70�i0�����qI3�j?B�i�Q~L՞����fIf�S��'&��չ�	��Feq�t>�E�Fw�K���a�P>���|��#c$���wY�+5U���^�=��Q��i�(��!���|�H����]�I��eԗ�\�L)k�+ƝwP���3����.����&f(ۏ��T�(P)]终}���\)hJ����
GX�:r�뎋�5�?^K�f2�͔���a���0���-�V��JBL_>�/\��8���g��y� �x���!e���Am��)jR'�e�J);Dq�h����;,M-LG�^��`8���:�m'�k�@B��|�+��$�9	fʳ�-���`X�l-��T���3�����3�1υ���;�|������.`=C�w��2둞ūc�u�w�n�9H�ʄ���Anri��p(k�,����O�ui���q�L2�I����G�
�n$���k_v �������Υ�;�}�0ܾ�l=e��"��;&؝�YJ'�R��FU�79l��r��ZF�os̻��樭�xU��y2�O(����g�M/s�ob*�$�E;�J���r����h���լ�b:�2�mk��Ik�;�ך��$wvo� @'��P��mv��v��|�3-��S�4�s��ȅ�̃�� ���2ߧU�\'C��ʼ�H��S���Gf���VƆB�m3Tp��1�G�گ����}����A��r1SFe/��Z����QϹ�$��RY�|��$*8f�D��d=[rî�������m��W2>5���k�y���˫ذ�x�c�]�4����~�,��R~7b`-���{_�mm��G�JѮ��sY�W%O�*���K���H_�ۺ��!_
�n^���ߓ�/`��f�.v��ˉ?����C�3-Yѣ�r��u�/�����)L�Ԟ-;ݦ�������o�&���Ndq[Ā��J9�7q�򎴒��~8l�T���ҍ]E�H���9����c  0��-=�᪕j��C<�>R�-�?��Lw� 2Z���U6�6h�uG�9��������م�|N��'� �PQ��ɍyo��H�b����`%�����J������I��
Gb\�.�uD�y>��EN��r�S�R��}�-]�[>!O#�U�W��6��A�S�Q�Ky��H��09<�pd����'�NF�i�p&�7��R|���8�w�9���/`���<���*�ߋ4�-�
ۂi�|�W���J��Gu�>�8�L7^��s�	+��O��Đ�E缣y�,�ܘE����<�~�k�n���� �Ţ�@�׀G����i�5�R$QL�S���� �5�a\��]h�8�9-�����J���)Dǆ��I�dH��wՂ��Jo�}K���E�2����7$]d\��1E�R���p,�;�M�6	�˼P�K�w�Wȿ����C���r�(F���c�j�=�?Ym���}*�����2��W��\ R1���	z6���3��|�л�4�G�ؽ�����Z]b�%W��gΨ�,�ۮ3�Q{�մN�7��5�1	�������X�0��m�<�����n�" Y��?�!�m���ж����@f�e;�G�(��,���� m���k0���T��A�9����h+OY5���l	�:�{�yVV
x�dÞ��>Z��,�������~��V�Q2e5w��2IZ|��iC8��g!V��o����@���nW���3�J�%*��h�;�]3���e]��\�N0?]��_a�ވ0[��N�6�[�9:j ����F���3Ds}��#>{�vdn��H���!��:a�cٯw����d�T���+��iH�/6�:�1L7	��Xm�kw���c�����9�W��!����0�Q��8ZN��"~���[#� <���5d��H2��5�='�z�3�m<�7�S�a����՚�f�C�4؝ÄV��ө`�"}�{cW �>o����ks��o�G�
v���D�e�K���}>ꗥ&�Oؙ�\n��2��	&��W7���3�׆ 

�L�KV��I�I�{!B>�1��I�]��h��m-��(WKw<d��!��l꤫�rNI�����1R+E�T%�P�!i=�Aɟ�%z�:���^�0&)���4:|��d�5��9c�W�၌D�65���1|�B3���3%y%d����O��"�BTD��)W��U�����{-��Ɋ�nv�o)��=�x����ORx(�<&�+�F�!�
w $�=w!� $-b܆���C���/>UT����poH��'�G$����t���7�2�"�8�c�Fl���7M���)d���V������͔�<�@+�ŉ�W�:A��%N�]&V�8�v[�������$]M�� ��F�Vu��޲�����3��c�D��A�Vat
}=Oܲ���fߨ�,rFl*��E��PV��蝔�V������c��A�7m��þ�b�yx�v��`�ꅤ�be[�:��C�f��Mr9���jS���'|�&H�(S�f~'���ޢ�$壈m8�����E�A�!I��hlA뻠��a�K+���u�b&�� }>H�\9�r؟ˋ4�9C�9��z]ї��C����>��0��U.Ϩ4R7�]�ѿ�I>\�;
�/4�4N�Y�ʽ�M��$9���D��ٰǪ��q@&c�(|]��l>��ua�F���
���$�V[��cX�Y�.���&T�7���=���QAm��֗��3M�X��;�^�������n�����������y6�[i/	���W��u-��c��E�6�Gƍ��B�2M�"y-z0���Z9���}�e�S���d.ŀ�A�JrAG+�ƈ����7qfW�Y<6+�l��֟�9��(���N� ��=�5�N4�J�؀����B����<~�y^� }!��ǡ8��e���{�|��˻�Q�M��N'L�/�
~n-�͎����}mc9K�YeZb��c���7([]we�9D[���������"=?`�Q�-��y�f}}R`9-�La�i�@�	�9 ��MP
��SW�ʞ�ۭx'vN�.�\$���T��F��#����@e�D/V�2'�~���i�J�%�v���ܻv�ɼ����T`b���,��f�w�nt������-�ݐ�:��\ME��v�q�io@\lҍ���z�{�.yxl�Y�8�*]����DR���o*��.?�a�ab�/�g>x��?-��"�.��S,Q��[ҹ����ֶ�^;s��`�q�eUS��VZ��4ګr���^0.� ��Ai��ޤ5D��� h|�Dќ�A�wm�as��Jʄ��.A�^f5�Ebb�qbJc`�8� ~w��=��d�}G���+5I�sa�49ڭKyq&�7�wW,�p��ON���G��+8�0U�&=m!������크��2EV#�� O�C'
�^�����1�˒@��/
c�(=��V[¹"�cx�Fh�hF�|�%�1�"�E��>��o�4�v�J/Z��`��f�	���Dn+l��^-By��^E~\_E�֮&�g��P��.��apP��W��|"1��������~i;3����/������9�q�$�;��
���x̸�����sF���<�D��{��d�F�w΋�s���Ǟ�l��Ұbx�څ�u�u���&���IГz�S�;�d���l�|c4|mϪM��?Ҳ{� �D'��.�� C��#�m��Ѫ>�^�7�#埕.&�`al�0�e�:�P��2�X&z+e�	2���%)�s�p>ѩ�CJ���k?��B��'���0���y[�`Ϊ� ՕF�z\I�9�0d���.7�E�i�Ӧ��2�m�s*�Ѐ�?)�%X_�`�>��oZ}ʮ���Lb��W��/�kX��)e$xڙ��@��pLܦ>�10��RaD��F+�J����6�M��X ^Im�Fl]*_�>��hC3n/*֎�R-��u�o�cq�z�7��ꦙ4����'�4��4B`���R]�݆B>^3�����ר�#��	��º�D@Y�;��2�ՂK���"��.��³s,��L�6�։������L�P�w��\C�L]�t�w�UK�֯
�Z�j�( 4sA�\����Zxݳ:x���K���[8��;��pA�ѭ�^���H�����f�z!���JW��x�p�1�uc��-#�nV�I3y�S<��<!>�� �r,w�4�9ǟ�q3�,8�˙Ռ��0 9,��hB�UR��d9(&5�Z����V"-��7"�B�	��`�����t�-��*!��VP���!��M��ߺ�Y��'zKc�q�L�S���z�jf����/D�Zěl�?c:7�ݛx ��!�W5f�$�)hՎ&��\�oUד���^Q�~&���>���.DL�K�f����M�yI���_�Q���#}��g��h�+� }1C��a�VR-����������@���bK?��P���c�5�1"V��73>K>lO��]TBm���)u���v����T�ēzV�:�~�:��[�Δ���Z�n��#StR�OmΕ2�Hk�Xצ�Va%�񗢀X��$h�}�� ���dԯ(TD$c#*�hv&D�ܯ}�ق�= [�t}zwE�Ol��|҂Ǣ/��#��<45�r=�FW�6_�b�wg����4i�m��^ Y�
��R��0�������4�~.�
}��F��@���H�6��lK.u.r��E`*H�G-�4�JTS���6L
���ww(~w#ۏS�ȶ_��B]^�܋Wk�*kn��	eQCk���523�Dq�]Y�Z�&��.e93�)1�8y�,y�����H�����ɹ������O��)�gb����o�叭��i�>FK��
J�8��T�e�������V� \�O�7"�l����.o�?�9Z�~n� l~��m���$�l�����ܶ(�?���p�b����ş�18�c�$V��S��MQ_Y3i���QB�.�`Kl��mm㎔��)@�&`$��Ǎ�^�p6�zu���#�>���������R�E�y�K@-�I��+��;����&��+�moR�:3�!M�����Jb��������R��@>�>����OtvH�_�]�_��i�o����Pt��aFB*�@�w�E��U���A�oX�o�Ʀ��Kиd2��K+GJlj�����lD�i����Sv� '����������j&�5��Y�H������T���S�rn�UѾf��fE�2��;��
��h�@Ϡ<�x��Ac�PCLn�H���ʏJi�Bo|ﰭW�b"���wf�6��ݷCvh�f�z���/(�t�M�`$'�A���ڇ#�ͤ�� �h�&8ؚ#�D��t$�&�2�Ä�ev�?v���G|y��׹��K�|�Z1�,v4��h�w�st.p~�Wu��`���9 �
�wώ/��ɷtP;�aF����j���
(��Q|������`��n��l@{3{t���wrΤC��9�X��ߞ����Ê7�c3���+��/�l�ç��j�;�5�"��=��]��~�9��c	��^��Y�l*�1�>�dC���}�I:�z}vk��˰B��RF�ԝ�,�m�'/u�/5D��8�&,V-9�uv��a�Hg�����{��s��Q��	��M7�п
oyo���E�f��jUc���"�	�d�5�<h;�
�WK��/8�!
���s{���bt�w��t���ǥ'h��)Y�$՞���F�2��@�|)�y�ǖ�3��}Ԫ��lb���S�O��r`��bO���Xz�b��"7)x�D)�|����W�kǥi���w4�qk��B�W"�A��^f��b���l���'ӓ�P�3<x�1����~��.����$-+b>ɝ���M�U�}qRnE�ω�H&�IT���+����@�7�F�@O�yU*��b���o ���y�3�rL�	@����!�V_3)Za�Ơ@R�,���9Փ������ss��P���<�jL3�=�d1�����^�0��}q�
������N�(��琢�3���B�"��ά���r�2�� K7C��6�U��)O�1Q�U+���!�'��Z�����s�@��W�>߸V�r����ԍ� ��\�����!�*5��,$9s���]��?��T��폴jyL����l. ae�7�s�tc�;y�����1�W�5����a�(��v{���#T-�+H�~w�YGۘ�׈�y7"�}�ek$�(�i�y�_h�Y��8W�1�$�DX!{|�Z6�T_����]�>N�/^�'!�
���Jϖ�{�U�T��=��A������zf]&a����p|vc��6�1(J=&�M�n}���kqF"�����y+3lD7y�*�5��)�-_���U|(�2ZVO���7N_���q�g_L�����x[^e�&�6��G�G1)�ܵo�ie�ß�ɓG��N��A���6Շ�:i�f���WH۲.\DY�K~x� C���`d-�e�ڻ��� �ur��h_Ԕo�[�υ����Ö�;K�=u�`��_M���p�̟�vޜ�`�'i�at����ju����(�C������<�?]��kD�e��ooz��I$e���F:����\f�P	��&�J{%�ޛ��>�\���vM,"�"\~&�L��.0�]K��Cd����}���<L49}����S�|�lA��F��HZ�$2��Bb�`(g;|�d�߷A4���@nQ��cX�>6�%��y����R�.0lU�
��P��?��
��r^�r|�ݙ��z�5�Zn����"�7%�|���_���mXa� �ہ�֍��(��U�R���;��ɺ?��0��@Sݻ��[�8��^1O8K�I��1�˴�-�h�4H��0.��9�"�ޣ�н('?f��p�2��O�uE��(DSg`L�@ ����hD𫡬L'�����$���[�����)�9+,�0:ž�L�8=02S:'$x��Y�б�Ǩ�'1��q+�:<(��o���<;�9��*a.Vx�>]�g��N�u��
 ױ�_�ПR9;�>�{%h��:� pR���`,T0;��P��u11?xô��t1MFSx��REh��S�53��ǲ����"^Y�[
�F�"�]��i�#�����Q  c��-����D
r?�pہ�qNp�hA�-�]��'.7����゠A�Z�sL #�]�$�:���Y�c�ԭ^+�*��=|]&f��ZB�HnG��A6;yfN��ϣu����-��CD�y���]r�!��n�e�ݘ�4��ev�%������T(��R��B�B�֖�`��.ał�Yh���fY�YǶ(�(��&��NiO�02����l�`��x����/�m#Ɩ=Yq|K�j�ڤ�Q#>�NՐ܃f:��2J�U�Wv���P�}2���o�9e�[�Z�s�vV��Ȫ�b�V+Բ)���J.I�sM�k��
�Yԙ ����A��0|;�̇�mw0����X��-����p�2TB��Ax�y�/�G�vè��J��zD�H��JK�2�s���'M�"t���|j�m��#��]
���x���_��14�K]W��^y,�ԖGq����xo}�!��(�ݐ�0i� +k��j��7[U�@ u���4���L&�Ɏ)kT�/=5ݯ�2E�{����:_:u���{Y�f>xU|{�$����z��P6�u�} ��>*�r�P�ki㲨���^��-t��5�v�Ep����]1��L�Ej��O����{n�qچ	�`���l�ى�>�)��@:����Y��h�$I�AX{X�lBb���R�[s7�xm��J	�s�
B�����I(C�������6z �"4�(�Hd�髿���?\�8���>�sUvI�c'#sr;'^I�1>z�x��V��P�/�w1��z��+���nSA�~}�������NzVLh_7�LxN�?Ф	>�8l��$h�]�+�*}Y��75)_a�7��
g4������E6����xJ���/��;��*��_YR��?���n�-U���h��:ja�G����3���d��M|T�G�[j��I��1�2<�J(P���I�a�$�DB
�@ɖ̂���y�AYlV@W��ȔEzVh�0� �\C����-`�Ut��T����[�wC��~=��3�Aaq*���|	��m^�ҥG�+*N��Y�f�Up�S�TI��0)�9m�,`�*� U��ƿ�sp��i0�����'����vH`�miŸ�Pdh, �x��2B��������Y���(>|�&`|ڎ�JO�F������T�.�7(���u3��g��H�:Qk�����Z' T6Һ�i�,N0
�:A�MI^rȸ�t&F^cIк�\+���T���Rs�L�Z@QE�ߎ�ɿ�tFP� ����%��1�8�;"�0���uQjq�Zx�2��ٻ�$�a�vK�GsMV�:qVf*~���2�Z��`%�q�`�7�eF"�������#ʟTZ-3�i^9���bm�m�2�0�h(�G.�a&�Z�d�5/�K�"�v���Mh��('��̲�������$d�uVI��p�5|��s1��;�����^RRK���F�b4��,m֓ӟ�����<�n#�.� �Q�I,�_��ף�
k��!����n�{����/P�̬s7=��8��*u�� ��B��aA9%v΍��qYXJ��W�� �����	���O ���j�,W
��s���i\��0xk0N&�����q[��?. �C�)3���[�ւ�5]d�rm@#�s�Z��[{5�i[���$҅N٦�����U���N,����`��N½V�r���Q�1��H��,��zA���`ǋL��{�8�Dƻc�"w�uk�gQ}��(�ƣr&�k4m�./�f��i��d82�p�F��Uc`}��c��9���d�k��8�=a��5����t�c���;�Q�I�b$A�t�x�8�D�}�y���V�3�Dƈ�[��fD%ݶ.[� ]��`x��K�Ag�
��򶼄M�=��{�;�K���}��Af��RI@�]����@��>����|T����%BY5��W��p�݊~"��	V���_� wL�kI�L�C5������&�|:��qKwͽ��w�3��X�1�#�mQo-f�m�r�17����L8O�w<���*�H���f\H=v !�\�di�.���byѳ�*��;�� -�eV"WcvE@����|��N6�5��rk��(ZOq�Ud��S�ߵE���e�ӊ����n����j������[��W:�˞�g�3�4xPMzz�_D����.�:�y��3�����!�`Nʍu��A�J����ە�����_���3ޞL&m��w�b��\0�����|p��pNX	�PZ3�^�a5S�K�!��ַ K����� ��`��������!ǒ�z`������s��	rn�7�y-�1�K��q5�#`NLvJ�/�zfam��� �½�"�7Fx�h��'����rDZU��h�5o���U"����f�%��0��xz���F� ���Ե�h_��f�Pu>[�ˇl����-X�f�g{�$U�b-<��e?j�&�|-F�<6��Ӓ+��H���e�8��@�G΄L���h��T=�Rk��єg���3���g��HUY�q�6pf�udp����@�z�mg�(ޫ�M��ta���UI��Vj��Hh�/����9d+ϐ��-�U`��G��󦒹i��o/3���[J�ߘ�ŒnrL�@�eoK<l��U/	����X���<������R���GBTA���B���u��Q=�.���f����R���5]�k�ק��\��z�"���*9U'j+*m�����
O2��������/kH7�fA�ᲈxx1��~J���ȞƤU�/^R����=���//^�;����Z�D_�L ���������?&�7����0��:b3�<=��nȻ�Тy�^xG?��,��Sp��'�ݜ�a���L��D|��V&$A�w�=�({�`���-j�CĦ�w������F��Z����4A`~����)j��'�ƹ*%���T����X_�v�*kKT5G}�U��wp�r�;�fE�Q������Ӿk��gN����UJk�8Co��g)j��r��Q���ߓ6 ��Ob,u�`�	��Qs �DTS-���o��)VH~!$��m&L�����E���(�}�!��$�'0��oŨn�V.�|JHe����@��J�qSc�P譭�3��J�ԗ��ev���B��(f	T[�������$��rL8~LbN�d1�Wf��us��A��Ә���n'i�[��J-Ϫѹ,�8��eN Eߥ��.N �9e	ڧ�L��r��Q*�r+s"���u���1�uV��C!Y�l��N���׌���6�B��m^��q���� ���S2�	��p1:�mWY��������wJ��2]��Y|�NY�"�n1dt?�s�����纥��f�:��i��?���%��%��r�;Y�a�}��0��T�#H�-���@P���V��l��U�X��,B&�h�~�n�R��~����\8�w2�J�[�����"���P���@v;v?��8	*�{�N��2��J~=��(�?�4��~�U�w���D�0�ko�m5 q/�) h��`g�]B@�콥.�%�I�<�{	�a�C�C�li3���X��
� �ŕ�.'ևh�)[C�$�z|���1�oͅ�݋.�Dvek�d�t�@	٠0"�1t�
�h�B��WB�F�e�+��e�������&�Dj�H�H�"���&��r���wG��?�z�ц�l���^C��M`[Sp��X?�3 Tc�u�~y$뜋�&�g�p�0�I���kL�2K[���̼:��=5׼O��w�ޭB�a �._΃)[�6Ef��+� �:��^�I��zS���=?x"j��N=Q��.���~ g��J{�au1�p���������"&8��i<�|]P)Or������R�-��&��»�c\0(Z1r �b�9m�tP�餒x��+��Fje��xQ�#I=���T5�}}��D8c=g�v	��T|�W7�a�CU �ufPW����������q6��TkY2�&~=$e��^P,����&)s���}���i�ơ6�(�%9*�$�t���wu��!�	���'E%�?�LaN˚�?Ľ�P%�^
&�ʓ�"uD̲�U�3�Ȇ�G���V+4�"�i=B������$�����O���d�%��C��F��KMx���
�1s��P Z�p�'���AN�O�{�/�L�E�h���=�а��������-�vU9q^���ÇNu���U��V�w���P5�E����S�TӉg�85���'6�ŵG�xܢ���Ƹ�5���A rX���ss�3xJbE��I^�5�A*�/��%5Z������-'z���ь��Y-�ۜ�e�p�"ۅB|Β���m�Y�rm�l��'�S��e���ZUs���x��[>bH�},���":�?!?(�b
c(��gu���;���4&g"]�߆ *g���A$�(�ܡԱ31¶�K8Z5����Mi����s<c��|˙e�T���`2�2r���A*�k��s��Va�/�aq�J^���4\y�~'N��S�w�
f�eF���@McBp��-���Жm�F�֬�8lCn���0�4�U��g��m��ܺ�-$kַ������p���@�������Ͱ��_O9�i�������D�#����)	W2��o�����.˗_>��TUʗ�_���8� n��iCנ�FG�P�x-�6_�q(�(���ֺ�h��[*Z5j��7%b*�Ϫ�02����Խ����g��,+)pB`��lA̔���w՞ٵ9U���^�bZ���f�TcEO.�^�3�n�͒�V�=V�A��#�Kq��O�N�B���;x,�83\籁�Y��[�@�h!���_��+4�R+��� �|7�hJR����Z�w����Dm+?����p�y{eN���~�߅\�d\����R���q��ѫh4�� ����)OfP)+ �2Ŋ����Z{ހ��$�E�i^N��'IU��X��m������͊��/IƲ�L~��p��ȥ����|{x��į������ ���P����i�šW�<��Q��UF�P��!�I���Ҧ�l@�%�~ka���,V��5�@z���B |a�l(d�����
fSn^��8N�'�������r�Хڋ  �[�'.xx1�?�;��5���&Xs#����M�@l����3`_�HmH�b\��I"�|��������^[&WLP����<�*HⰕcۡ9��FWZ=����[�F��0������F�s���½�U�h~���&�?T�Ab�n�ya�;�pY��{�sC�G>6!jD�Ӆ��[]KG��T��T���qc,Xe�d���LQ��VP��.-���?���}�e�W��_�'�ǘs/x��xjc��o�5oʭ\��?�N C�ǖ�$;k���D#q�}gv��CX��x����Pdiv��	���/Bw��4
\����� c÷��J���� }&��,M�
�����Vt�u�G�m��g7܏�gX�eƐ��s(ENi�f����k]!f�A91d-4�|�fߖ�{1����:m۾"�2��҃��Á�����o%w�8��4���y-���O۰룑ɲ����s<�T���c8�JLϙ���2�fT�!��5���W)F)xD;w��P�"�Ք��؀fC�'#� ~@��eZ����So�~� w�����υ��VCW�~��S����6 �W\];ra��F� ��(�e~���Y�������L���	p�%aK$mT�\��@2�yLٛ��Qu���GӍ�Z���W��������e���̀�1c������h�ř������wsZ��f���R�y���>��(��5�Q��E��>FU�9g�f�:��V���]�^,�T�ck 5�~��O�$e�{#{6{��A��L�e���|���D`��K'_�JUv5+�-X����;Ɔ�
��<���x�5�[w�i+�q<�T�{��c�R���b�9�iB�	�\�/�;~��NJ�����+��?p�!�5amb�Py��������VZ�f�o�̴�암4$W���]�����>�7!^ԒH�p��e����5A+��L?
yK5jA72����]`����p�[k���pq�&��s��[-��N������5s��X�4H� �n��Dc�=,�;{�#�S�����,@ǅ����VM�ь�NI�������9X6�fǚt�57Kö�،Մ�2�	�O����R��e�E�#k< ���';�mH5V���½F�� c1�UZ� �Ł��#jI�4`+V9X����	���	�n/��n�I���m��
,��|���v�Rg����Q�3G��	��������d�x{�HXd�,�Mx��d��%Pf�ܞ�5��n�D#�X�'�h �s� b�3�b�h��aq 	�?qs��I@�ن�#����.nFx7ehy��Y账{c<7$%m��>�����-~Dg!{ӉExr���NwEBk�}F��Զ��8 ;�!�;/ns^^|�cX���ѣ>�"�����=�%�nr�N�S��н��@Bc����1nZx~�_��w���ʯ��
���Azoy�z�*��nb?����K��E�k�� ��5�R���T��E)�/l��|�5X�Q�6>�����a��m����Q�sʢ}�..&��!
V\d/��~/ex���D!m\�W$��ŦB��r�,ϴE���4�4
x��ZAmd��<9�6���?t��;n��[A��'S�좗8�%�����\ʽEם��q��g�A�ku#9�51~}��l�	��R�9��{ Y��B�ݵ�OC��EmN�Q9NqԵ�|X@9	�CߟE�!u�5),}�j��I�Ўf�^�B�c8�r`�ҹ
w8@�)k������o�*��s�+����8�[q0G��Q��
i����� 8b �N="V�y�P�c���5��]� ����m���-<��E�Q�@�z��`��HLpL�(��2A�A�ӱ<-#(!y�c��;CqP��� ��x� ���g����SC�_�,���'�n���]�S
���r|@eʆ�)��I�>��6�9�U�[rN�*�R|�Q�ݕ���Y��rS���"���.��6y\8yM���N�a�kg�O�C��#�� Z���d�X��
AW{_�!ToY�1�M�&�;�䩐�"-(Y�W�$��b3Ç��an�t.��H�����%��-��=��z�]�3�sbt\��J�l�o'�Zs��y�DE�S�;���d�_1�'���u1�^=?дjX㺷���}Z��8W`g�2oL�$��:8�̢��nV��p����|t谧v4CӄH7;׉���ф$ΙQ�#}S�i�)o^����9�P:�L)͈�+����U	��.�hg{�+�[�~m)����('%�X��c ב|䉏):�5�QT�h���Z|U�ip���(D��Di���>�#��*�|�HZK:v��ޖ(�J5��u!����'߄��4g�'�J+I������%�@��F�݁�xB���}�O{Nr�aT���m2��l}r������郷����2��Sa��Z�FXt���r�1N�_~;*7��5��"Cj��"�--[�k����S�	ł/&���B>����;ЎXC�	�[������ޣ���{;��|Z뎮X.�o (iG���Ή����j�ť�'���w�q����3��U�>!���0�Y-���Imf�b-�
�{�hru}nA�i_�e��K5éƿ@�YKxx�Hf�z)�ixN�F\O�CY��;pi�yK�������R��U��#��} #�I�D豱j"���y�	©jkz�s^FO&�:[�<��.c1����G��9d�zw�A? ^-]�*�TOr�O0�B9O��*0���e����`����I�Y��=���(�R�hJ��y!5��j���*c�m���Ce����^Ŷ2����y��â�|w�	��Se�
4� 2�r.cq9���
��3#�Oq�My�X�L�uKA��9v��9X���=�h6���� ��L��d��w�l��-P}bB��bZ8!�Q���'M��>�;���ݻ݅6��QD��.]�G��z�M�H0�,������ WD�@�T���!$����|�J�:ة���6C�Ҏ=ٳ�+�P3�dMn
\�*����Ҝ$��PIB� ]�">d6E��O/韤v;g���YM���I��I�L[�d�u_��J��0԰��U`�z'��j6�����/4}G_�y���6����八�ڿ���gd�ϛ��Bhk�A�8	w�[�﵄}ӗ8��j���[.��F��]v3�r���7:k:?��#O=�}�k����H�7�r�
o�:3FA[��)�������jX��[֢y���І_��������/�h���m�$�x�j4L����q/�`�\~8]��t.G�;Ĵ�FK�si�Vը��nZ;�En��]����r�]��ot�ڲ�r��-�K��h���"�[�E���)�m�/2��	�Ks�;�-�A�E���>���LnQ�>����#�������۩�;jP�� <,Z�ʫԳR:
���zKWߎ�7T'��r&֞���X��4Aa����)G#Ьj"�]iI�-����UE��z U��洪��ߛ%��МD���JZ���5gJ��Q�8�aJˬ\T��i�3��\���j�ԍ��x�c��_�C�����jj�cs�#S��(���������>n���kR���z�|�$����	Ѭl�|�A��9W��΂��(tf��(��g��?�#�Z������/�~�si�m�$C��?Dx�v�M ȧ��#G/dl���9٥*S�0+�w�� L�
�L�_��U�I ] ��M3[ǟԯ�>"�M �n�n�ϫ�����<ƛ��Ӻ���}k�F"�һ��䪣:l����(RF�t�k���~*T=�z� �>�Ymo���r��.���y����.p�1z��b��yS�h��:><��@�3������Ú���}���v��X�P�B-�"<�g��*�*gz��u$�J]��2%��&�L꼶�'���W�ҁ��z�z��eSԡ�xb�w�vx��m�ӿ���%+����4!*��L1���YM�#+�qCw��P�%n-��I�e�
����:k�y�E�&��=?Ju�䥙W$b>��:/\�.�m���s���z/�E�̢r�u5�4Hۊ��~A�#�����/����eʪ�ȷb�B����Z��&��}�E�X	,2�Vq���Ѡi�Cn�X���&�\)�?}�7���=�ْS���k���	Z� ��'�o�qFtH��*RUs��g���
I,=���qMi.Y�0��3��KT?M�P��Մ�p�%+�@�ws~k�v]��<�Z�,��+H�m�XQ|��o_��e.Qt��z%����Z,�'�57C���jLҀv���^dB�K�2\lg.�z�|IG�r���d�]�[���G�!����F=m Ky��h��#v���#�3^}�c�<��o�A�r�ۏ>�=����N����W@��'Y���ǹ��/�#0P��b�X�<<R�?�!:���p�D�֖R~D)�(�_^͑BۺCG��]��nx1�u-��f��
����Ҟ���'G���SB,C2u���dp!c̣�x�$��*�tPK:$�*I��-v�CkFm���O�W5'���7���"�߮�����a�<����]ߑ��}�ۦ晓Ii��J�/��)FP"�޺gN�`��X�U��+�gl�R�i���o"�87�6��K��D�gEu��}i�46Y��c�k�y��(�qԕG=�8�{/j�����X�{~��[h�R(B8ȷq�"�m�'�)M����>4�,%}j��e]�О�)�(�K����(��X�?i0��Rxx�d]��
\ ����?��xć��V�l��Θ2t0۳:>����������Y�����$L�G�l������ȎZ	�uN�)�v" 6V,H]x�v�l�f�ꄗ{K%�z��*R�_u�.�k�d���/���������^��-��(�z-���{v�E�P�߫Qa����;W�B{ݸ�7G��u���ai�\B�[������^�+�kv-F�dY �S����>��'N8����7&���Pk��X�ƐJ��û�S��ݩp��C��\	�i����Bb��*�%���<��]zB�
���±�����=�`����\�O��@��Bڭ�H}''��!F��<E�|�n��Ԟ(��q�~be ʵ�Nh_��M%U19Q��E��׏���"���&3p�>��c
��Bo!���
�d��T,�L�/��m4M(�<���u��KqmZ1n|���"�+�U`I���qy�����rhu��D�2l�b����pd3���Z�A������WX�a�
��n�^��zj&_�|��n%e=���}�a.Z���Zar��h�f0!84V8����G^�L�϶?�����+g������2C�	��	�V��.�FCQr�P˺�O���Ubc��YL�hֳ���X+Lb�s�H+����4�Ԋx:�ӻ�,�q�������#�p�ч#µ���"��.TP�ڶ�/zjn2j/���9ް��H�bSɰ%K>0J��t�~��,�f����P�]�?��`L�v!	��7%JrC#-��J@,J�N��*����O��kT�8񵑼D������ڃسpr�����ڀ!N���Y��[e�$�`�fU�h�3K�c���`����2r�Ho��iا�����Mk ���Ь���@���@��m�	�'$��Ӈ�:h�~�}Ղaѷ��A�N���a������43�&�����.��q�#��5���n��&���H
QdB���GE��%��P���z��u~C���v=#���,: Ъ4����'rl[p�c��ߗ�E��0����0�^k��1�Vx��v��K��g�>/��h5��a���Q��}0/ <�#>��;��`dC���w�p�B�]Lr����ܬ�R��� dj��M��z+��.���Ϸq�ፎ}v��w(��>V@��[j%FT���mG�1q2�쇯��G�6nb��y�BI��b�:�	�$qLY�;���Ove����d���S8e�h!hc���N���&8�./��Ub=,��^��ӧ-1�̥*�⟭�,��^*�[<���G�>u(�L�o�����P>�sg�˰XW�IH4��ff�>T�,��:1�Hԝ���UIi�+���X��@.�� ��C6�Ӌ�r�a�.`���J�
��;4��:)6@Q�l�C=���ޜ�<�ײw5+���XF�r7��
�K845
 ��BE�����eÃG�]R������-aL�Y,o`J�RS;�k����A[�7�Z;�1d_��J���E�u�f���j�x�F�A���M+�3����v��'o�+wb�R�7>r�q��8��E�DLk\���	�{�uvL�!I��s20?��<�I��Wf�Q��X����^(�4~/�W;E�����t�\MKDQ���2���(�ntl���nwm3[���{�
_G�`hŜe|̱���C��*��g�����g���ܽ�!p��C��ӑ���'d�|(�h�mK�ܽ0���@˿����/[l.��*%�}�Pj�����n�b��32Si<�����^�[3����Yc�=Y*�`���"-�������˘P����k]�I��8��^�����F"تeDq����gI^�a7�hXb �#��)ɛR{���_����۬ːޞ������3"	�0�#��z=�>������j`w�]�-]O^Tr���e�b	�p�T��243�KuX�	���R���~@[�.Җ:^oK�M�ۅ�}7W�4�i�~p��9�P؁��Ā���[�k�w�чP�A��I�����p��y��45@�,/j�ĥ?b�L��)g��q���$v=�_���﷔��*g�;$���v
}�Y(^ 	��\}ȍ�?@�P�7B��s�L�c1�C�9��D�1�,�t���#�;>���>w��f�f^S��hJpKd�m��P.	���޻cCf��n'�M������Q���mذ6?��1��/�� ��^���wH˺��>M-�$�j�{m��"T����8l���TQ7>l�2�ܕ���$��2S��A��q_�� i��b�b�z�!���ب�B�Hℯ���I���H9w?�� 8�4�< �|]Kȭ-3�+���=��i)�ى[�H�T����L�i�2�jTV���X�Q�I��7�\�4������]�����qW�ǛV�οK�(��?#j%4�NSV.lx�^�_9T�g�}s>@��$�<A�y�l��5p�Ώ����|��a��q?1�ϕ�����J��w��?婎��/#���1������|�2���0�m�Omo�{Q��y��~���<��*����>����lײ��6Խ�#�'�D�£��v�e9i��!LW���6?�ރ�cr�r&���J����+s�<�'�������BdV�A�:cG6�w����	/��~�Q��Jzz�}^ p �y��`��q���8��gU���~߮8m���|g?X���'�<����?�m���??߆�.����eQ�C�f����ɺ�xC2�w�p�byEu��0;�f����Y���4��ޛw'K�us�?	˲���!?��P���:�l�r�]��~:��Fвgm�����%P/�� ����	`��b����ۥ�"�2�8���db\S�A�Jv��?.J�YU��3�^��ʥ�$�C[֑<	K���D
I�iݍ��FWL�����z����V0K%�a���n0Pj����6N.
�e��cD��Y�#D�/9o�[�^�˜�����۬PfYj���%���ˇޙ����"Y=���Ը5Z�d`�ٛ��)r
�ZB��/�Ǚ�#Q�.���GI��l���m?W�J������rs�n%���{��u"-�DM�]�89«��B���P�wWU��x��MB��\V���x���on�o���`yv�i�h�]���uti~F��i����7��mZJ'�GR(f�f��B�ZL'�S|ؖC�H
�5�-V�;���C���))|L�'^}p���Ͽ��n�2oO��N��e�	�p|���������m��T��^���e�7!O�;B���DqX���S|�b�2^k��ǵo����fñ�o��6h�G���k�1�b��g�]��;��1�z 5S:�D�GR�ݒ�|A�T��C��	Z4	��n|i���=ϕ���7FIM�T��7����9��moLXn ^B���	yx�pv�Z���OQK�a�S��ܰ z��r�՛��ʹ��L���c��\��y�A{����|�"٫cT3Q���c�y�voך����;0پTsS/;�I������ݭ8�<�Nh�v �Vް rBIy�K���A���d���3�'����,�9�WEh$羅kI�`������ v֙ |�U�<8z'���ϖy!�@-�#�ՙ���d�����	���]!th�,rU4���a�#KD2�M;�حf5�"��s��a��Kbz����H�d�5@Al�9��XͷՒ��̵'7��+{9�G �H7�p�ZW�+&a�L�j��g�������8�4&@�f�B�5�1v�?�/,�~.*�!i,� ��5��)��!��_�Jm�t��OI�^΀��-�$����hl���,t�d�\���L6�e��)T�sQ�,ř�l���b�MU���t��!F�p����M���35QQ�4�����,���SQ�����O��N�o8���ї�|��W:1Լԟ�g��-l(���A�+�J��c�t�Ҍ�:�a���v�/���LM�c�n����m�q>�d�S�<""��d�l�H7�⵳�\���3@󺏬.}�?|t0��r�d�+!v�3*��N)4o�_���Ѻ��	�o:z⡪o� ��\�~E����qHITYI�q��^��l��1v#͕���t�t����K^z�C������m2��������4t�It=joҀ̏X����d�*Ҋ~�v����P�@���^��"�ȫZ��nΐ�yhr�~�Z�r �BU�a����_�HtH�=c��*"bT��V�\��y��$]0a��f��*�6@NRw�4t�����ͳ�m�;�i�,��:��̯�OM�K��s�_�z�^3	D�"����J��Ci�����3I���|�3ŵ_8�N�|�p�̧��5����.����$>�:]~�2��������VNmʤ�ÙxW����$�&=7ϔq�A�V��+s��U��mmKjw��<���גBYd�b ����2�DH"ό�Bg����U�jV�_Bf�	��K�]��.�e�e���X��؂E����XUX��A�����A�t]���� ��' !&�! �1M{1Q���H��o�A�H3���-�#�ߛ�0�F�kc`*^b�\W��{�*���L������D�����#s3�k�y���f)��#>5�<�j��(��0�<f����1��n�VDVt�J���%��Rk�,��*�{ [R��hp�K*y�:t
�������F?�!'( Տsl���U����r^�i@Ħ�dL!���{��A�,���Pd(��>�vk݃~j�p��O,���h;Q"SL�t��%���J��؇X�Q��U
���TCQFS�gW�u�i��
%T�)�U��ઐ��mь����ׂ5Z���w��=�96�ӭ�|}��V��p��?�F���R�I�B ��z���5�X�umLA8��ZN��+%Z<�;x�� ~怽���>)�p�/@��ۢ�ϸ"Tw�X����}r��6�	�SnM2~�c���[��b��C|�) 6f�S6̳��B�ڤh��ʧ����ķgd�կn���5����*�~)�/����7�C��M������R�ǋ�j/�3�n��_�֪��Tܚ2�ł�5M����b�m|_Ӿ��Y�����AK��!ō��E�yT��a{�.6���.�5~I���=}��Ǫ��ޖ7�l<c@�Z�~%*_���?��r��ÛD��s�B�-�DjnVk3��!�J�B����<�s��+V�B�>������z����/���=�xit:*�A~�poX�����!bx2)��S9�I�V�G{�7�.���YUϫ�7�j��8���� 9
}�<�O�9�E0���Q�"�'D|g��r�1���@a�LD��b&"�3���s�0i���f)o�M�GbꙉQ��Z��&r����ڱ5�z�x�w�n,˙�|�S�,>����&�~ˢY�PF0M>(���-����n�~��@�0`
�@�CHd>kRQ�=���U�/������E%0�VD�����6-6�� �Ʉ������խ�c{��O0S˵�W|7��Zz���Mw=2e�=�X���`�k)��d7
�l;�H�$��1��;l$���*���Lgk�r>��rtǒ8?5,�7��6�؀��K�\{7�9f��u;A��*�WrG�-ࠁ`�c��V.S/ȓ�p���S_�]��%G�m�E}[��.Ų����:����|8�Vr9�6�*À��&v�lg"�)R���u�뙹�s	��1��Sl��ћ$�L7��
����d[��s��1��-�Lj���Nԋl������jWD`�l:ax9��jr�g��'��E���n>�<@2�����]�3`�擗XR�R�P�+���V㷤@�{��ħT�wpi�����w�U�3h����J��1:����qX�����q��0v�#e �%�j�L�0�~z��/;��x�Ј�����JDDӅ��u�X@t��Z#�B�y��WO�l�O9�I��aY�(AkH�����3�I�}U�s�#�If|��2�1�DN�V�2c2v(9WmL�PM�М�r��5�e���������K�� �:���DV�S]��8�}
��3v��:t6M���6����N
}|bG�``T���.�� .EH�x���d)����ۚ?0��>q8��Ǽr]����H'�]��b�N���<�i���\�}���D�Z*�9[-I���Ebhݮ)3�M�_{VSX��i'���?�败�|�$,���I�ѨIۨ��sp'O�Kl"��zndX(�ǴW4��7�P�T��(/FP���+f�n���J�����V��,�� �_�$3��҂�K�	W��Y;�����E��Xſx�t�A��e�@E�����*�{I�p�+��c&F��j�
��1��
s	�!b����m�h���M���+O�_s�\M$��e���)S�*�:����Je���a"(s!!����o�;��K�SZXo�P�H��� ǉE���?�@G��&Q�QՁ�ϱ�گ��Pi]���^�+���~�q�S���p���ԫ��P2�T�+�h\�>��E��\�����0}n!.�� ]�]z#bF�p�ө��ܝ��~62J��ҏ����!���n� T��R�L8��*��5�8=i�p+W��C��-��I	��j�:�e�Z���9v�CWm�mP��`/�!�{���2�e�{�����OV~���L��g��o��:�φf�ӱ��o����fce>Z�,��?�e����T���J1hBk���a� p���r��KL&If!��H]�iK��㱑n�A�w1���S}=�0U�(�|���꼗V��V��~�&*g.�t���m��q���@�ӈ*~���o��rx�n�[�u�s�qSz��6�؅�u0�w+�� .��c�C�N5'
�#Zh
�&��nOl^�͗d^X�9S�8Ē40o�����gұH�ڤ|�U9p��/���tos_m���~����-
��@��X+�y����Kb�y��D�����7��yT%ס
� s��j9K��~Tyu�!]�a[d�����vlP�[k?�$�m�+���Y���R��L�����/���B�����?����M{���7ީo�;�)��%��x�>��~<>�Y"bk[�v��9�aޟ|y���z�w��2��cǑ�}�f}�����,��F�z��z���)K`oh�&��}}
��6��y��ٳr�Zy�؟��S	Wi	�Эz��!?n��=�c���C��0;�;�^���Ǖ��گ�k�q�R�l�~ כ=RM������PL��Կ�(��O�cBȇ���G!iO��K�h�N�,�o,|s&& l��q��:�u*�u���[�vժ�O����	&.\}��5YC]���sPx��Ȁ����A(�d2���l�K��;��C13c�Ɛ
��Wn���Fb��ݜ�����i������f�1��,� @�V�+�㧴��8��8����x���z��B0c���`��;��#y�¤�z�y����9��VF*�
�x+|%�����O��V��ᢔj�RP�zty�K�=
���$6�� MX[@ҹ�,-�e8F�[0��ޮG)��a�K�ⷆ@+N�n.���CLx,���8�����=�]#������U�<�,L8bxS��A�Rko]��i����Oz��1�|���LB�MlHgE1@��?��Ƚ�M3�ZE&�r�d��,a�;��Na��?.��0�Ϝ��>��2xƀk��w
ە=�:!z��߂�)���o�"O���`ll*�8�E���7��9:�n�FT�/IΌ� � �V] U��]��\J�+X����d�G�=b �F]���J������)�1 �,9��/��U�\�'6�-�mq�:r�e?kq�#!9�d;0?ʘ��Y��Sږ5ГP0 ��xz�tT�~@�$��?'������M��	?�t���H�h��;�`���R-��8c�d�-GU���G�en�A>o�""��Es�Ӯ���ʍ2�5�ǯ�5�BhD��6FJ����^a	�_ʟY��&��9�����)��VwMh��W�
�lօ��%�;����/]"��V�ߍ��~�㉐-R�F�>�׆��	���lf�����:I_�?C��nE6{�B-L�u'B��.YW��z������q�{�0�PP��װK��#�5��u2�Z�P��жu���a�����M�1�p�t{�0�R�cL;��h�L�Q�Z��4��H�UhJ���p�P���)sz�[F�t����y�;���4�e��Q��	�@��&������B������q����k�Z�6��_���˕<�C]H7a{�ާ��0���5�)���?e�R�ɑ7b�;�VUD�
6���uŷ�C_J����6�U*{h��Nf�c�a�=@�C�ip=�����a}�LKK��`�� ����Tfj��֣pO�p- %�g<�-�~o,�+�Џ�T�2
|Z�EcR�eI���7�
ew�Ԗ����?�.��h(Dw�dR�}Q��/G�o�eq���CO�����2M�H�U���@����9�=�"2&��&"��\w��O���uJ�}2~��"bx,��x3�ٝ&��P������ƶ*�G徶n���'�8�{���c�Y�*�A�dK�s�v�+��|Q��E��ّ͢J��,����neVԥ�(<1�@#���?���.��[y�%F���E��p�?U�C��=��h�񮂯�T==�[$��)�)$�l=@�'�/��G$�y�	٣  �Ĥ`�`��� ى1�Ƨա��?�� V������	Z·y�G�{հә����P���6d&�6�F4�G��o�5��Zh�BOY���n�F�r�<�s�,��p�j}�2_俥 �'��ñ�
��M�8H���M>α�.�k������x�M)�h�E�clB+!ِ3�7S����<ª�+2��_YqZ�B��8$ m��f'g,�[���ҖMnq~O�ȫ�Q--=ҙ��Ʊ�?���`��$@����I����߁mL�4:gUݗ��v)�y�!�o�0� aF��� �݌����wf�E�*(�8�'���^oΌ�a\g�EKR�=��
ҪHi�)�By�*�ZgN1;i���g�$Z�\;�i�����բV�P���i�n��ZY@�7�а$�����"���3$�0���� J�=r̋u��N��C�5��h檍��"��һl�f�@9Ғ�${�^M����q����֟Q�O��^S���k)�4��P����ӈ#��@��:�;�vǣ��*"�+K�O^�����j�t�~���Cңm[�/9 ���g�֥˴��T�����#��}�-�
6������Ӝ	�p�i��c֔?��bd�g��Ot����S��Z��I��rΉt�S�DֈA�(;o�E�1Av�C���4>�"A^o�����Z�ڽr�#e�ɰ�.�4\�#Z����ɩl�͐��Ib�5��K&�V�7�IE"��gF��A��҆������.�v��-��R��1�,��%��d���!��ߋC*Ѣ^ %��q3r��NP*��6�ꛮ����u5�]]�=�I| C�>}��2��3����A$��TR�̞��e��~������;��o�F���@�3��0ܡ�N��"*B#N���ڏu�Z㰲�şQHb=PĨ����Bl1�������۲�.~|��ے��E�DƖ㔩˒��cqV虱��`���%�З����3�7����k��`�^�U}���������lOtcHh�S�5;s�VC�M���-`I�{�j���uc�=��DCH�H��������_�0$]0C���=��Z��{�[�۽>c�Ü���{�͟q��Ӷm��^�]ԏ�2�����JJ�v��i���V4IE\����?���xZ�$'�gQy�h���ι��8y���T+IfTxA���I020��t���a��s�7���Vj�ԧ��oǯ�,�s=Zq���x?D��C�,�r(�!ZΟy�i{����:�O�$�h�I�?�8��v�������>�5G̚�Pۥ������+|w����)ɗ�i
�f���qrV��U����G���6U��w˾d�@0hV�)8�q������:#��7~H?���4U|����GS���n̴���=B�S��Hņ�j���},URI$+��A��zvTu�f�]y��I����n0����ɫvJ�/��� �S��h݊��Z�JW��MAX��M=����	^�&vN|ס���)�u���� T7�d(����_�_?g�;�u;���� ;ە��/,������d��|QI�ޡ�.�o�(ԈHs�{/gq��ܼ�b�Z����=�h�ߞ��0*n�6�v����_����;-~9r�xs��K+�> ����:	���<v�f[+��R��]4g>��U��R�s��S�����R	�jitɠ!T0����s �<�=���8�U`�=�5��#���v�@��J���t�ц�u��^����<����))�,S��	�-@	 �)�@@R��z�>�t}��v��1����G��&�
���~2w;�u҇OLH`m5"��)�㱣RBcb�.���i�4�$&"X6l���(� ����ߎWX�}��AM�E��vMT.a�]�t -���I�s�f%��}lgN��ږ��:u� ���4.���+b9R�j�~1��������m��ָn�H��L`�
�]=GRuJ[���{����������	��J�L��F����m�%(�J�V�������84vm��ʹ{p"{�o�m_��Ni�����a6��>Q��A?Ӈ�1����\B�i�kV�/��H)�	��Y��$2ś��l��:��n�#v%a�����J�wml���xX�Qϐ/XXGv+'.�����$kD��%�
�w8.��
��WS�i�.R���+?����w�������: o�s)`�7��������"�͍t!��239F�I��!\ў��%Q�\��!p�^��է��$lݨ�Ne���G�M�D������4}Y����T�\��.ɏ�P�imV1}��|�2�3;�������
)�E�O�-�7�l�/m�tb��n�����T�T��Zձ.�ɶKFl�A=*A��%�GћU�p���1�����V��#"�~D�NΘ��]�^�X�F �5�^��]� *�V��	[��N����V��t*\O�@�[ߍCb��*�Ј����#$�_��J���Ş;j�ՔTrO�!�ێA����&��V3��"(��^�Y
^�<".'�^�C�,`�QMr}�}ܞ�O�2����_j��T#�G�ы�b�-W���}��� ,��k��<jqEl����z+|«-~�S�����@����J.�e���hE�cp��%E�� �q��=����U��k�kh�{I��×�m�(��f-��A��݆^�D��XV2�T-����cv��d���X�kx9jm�ݯ2�s<ģC�1�KP=5O��,~j.����c��t�Ȭ��&%w^�\��K���ǜ�)�|{('׷oO�9�(��f��{�J�����N~��(�T��q���)n!(�M�|�#9hI=+��3ɜ4Z�3]x�a_���$���Ĩ����K2[�Kl���3SJ#W:���!��7�G��6;0����1�^�C�T
\� P}��߂�*����aa1𗪃��p��q�qG��k�6�ZFݘ'ر�� W�f���S<���GJ�!�)�1��a��Ԙ��>U�=c���� ��3��d�H4mb��֬oj������R7u�n4!Z, ��b�s�L|yD�ʴ3� �7ퟢ>�8B3'�ޤ�����
`J`�M��N��+�����c�_]�����4@�2��;�K�����y�dT��F��V�|m���QmI�2��	�QG 媂����և6"��Hl��1*Y��*G�7��n����0�g�xR�zz��?��3e)VҋE�q�(���i�ML��mp���k��iF?���j��W�ϟq���e	�����k���O�8����+aE�?�;奞ᡁMw������K����E�����!Ze�K�� �L�f��\b�f�<��n`L�en_9�xc�R*�Ƈ�)^��L�]
�����
$�_�f�[F��>�#�P���؈�
��-�LWA@+�(��l���? ����[�� �J�Z;c�$q��n>ih�����dY4�����s,�6��b\�@��ĭ+��!����X�kD\���0#���
�+P�/���
ўa��.�A�vh�DǏ��c�{������I��Ln�kA�8Ã�}��{n�t�~���>_�<�[�̢i�#%��z��q�0��ޓ��R���!C��(��{�R0mfzt�Q�r�U�1�h.�x�������FAM��f���7t�F�`��*/�����Ъ�O��=7�UX�Ȇ+Ȣs�ʮ�T��z�@��OG��~,�v�r_�}5��H4^�����gZ��`̖���n�R#�Ǌzԛ|��q��Q<la�C��]�p�0� �W����<q�L�^h�kƁg?�W��������PY{X@���H�n[x�c&ȸ,�]K�l\8���9��07�Y���ɳ����Οv��̈I��H�}m�ю����2y�O"�e��d>l�:�J?D�9���Q�%��1-���Q6bQrU�A�n��9/��J���f���פFi�(�1QBV}y��N;��I�u�����k�06Ʉ�����SH?�jO�
�ٶ������I5��Y���Ƙphr���[���sV��ޔP��+"�qB��$6���a�&{�x�٥H��h�P��K3���M(^>�Z|�xu�"V~����04u��J���
���綅U�X�:��1���x��~b����5�����_S�Lל"�,�L
c�X)�7^I�ڕ�W���Pg1@l:���h��D�k��\�B�Ќ�f:�w�B��2��kz��eNGx-0��!+̍��9� ���L�����Z��c7T�H��pz|�/�A0>����(G��Q�%�
Y1ψ�*�o���U�e��������ǥ�#��ր�� 4>_�ޚu�A
�VF7q����s�r��F���؅����h����TDRc��Ӡ�ïzV|����yfl��ȍ�P����׶o�N��H1�ڀ���67��7��Z��ܯH�	f�]1�6Ar�]	ڦ��a��?nV���z�_;,��bM����C�I�{�"�0���<zu�h�mP�8�y�T�0x_�j���3ӣ���jZ1Sz��f:0P��҉Q�>�$�<���Ӊ���+2��IaaNf �2��k`G�Ћ̗L��Iu���a_[=�.����Sn 5ˉS�cd���Qp��={�l��bp�(x�a������V�/|�r����>t�/�o�;��*:'K�>��I���%)9Ò�8*����GP�����XN!�%����������",f�-MG���VL6��4�\XΜޚ!ǲ���Y�L��X��D��UX��j�ox��S�0�a;�)5(0�5:�-N�N����z�?v����r/{=�_�Ri�<w���w\?�<$�ߦ��_��Y���F��2����V�x��#���O�f��<�.��&�kCZ,|�a�+��,�7z+��#4ê�qЃ��́be�nS�>���'	][�ި_��\4���Q1r
�3�|pe���Г@,� w`#�4�#G��ZRD�lI������{�qp�^x��7�1�s_W�~�f)�������\��6�����N�	P3�H��y��?1Nm���f�pi,x���Y)#�S�Ko�����Y�7`������Cf7j�⇁u�;a�˹��)f��Է����s�#�Α�bD�9��O�Oɒ��K쮐̻���v��u�И$M0`��6�o�L�~�RA�H#5����F=E�tP�wܖR�e�C����w�<f�E�.�q��Vj^NuU�g˲��UC�L��f�ЯP�;&�.��a�.�e�h_�C��s������{�J��	ti����T"�/}�R� �!���M��V筮M�PY574<����$h
Ә��
~\�uԱ«��c]��	W�ٚ�eU�j�XE���+�;�Nbv���֛&S4Η���4b�_mh�h7:݇� � ���1q�z��e�ݮr�A�J.dh߭<��n�ըx�#pk��؟�r�i	?O��g��=����4�y����u�&9�����H�̗XT���ѯ1��S�0��#C�G�;*�`���Q��zG#�plK�"T�=h�
<q&uXcR�:�o��.x��0'@���ͪw���a(��]���y�I�Gs5���SZг����;�5\ݭ� �m{~��KU�VRDmke���~Jt)��9R���I�K�ʜv�6*bEw���ky@�tߨ�B}o��k9�2��)�4X���T__;�|�Q�� ;/�$�vF�+�g��0�i}�� ��������^�
BI���xe<Ku�����ԧ��
������ph�<��Ӑ&Uw~�6M7�����d��9���[l`������,?q�?��E�9i��$oO��D2:Q��)��2K�:?<; >��^ލc+��	�N��%�x��K�]+��\H��v�����y���KC��A�؆�
?����X�g2n�p��������9>rlGƪ�tv������,����WW��������V.�wW�e�*c�]��5��¬���qܱ�N�4FT��f\�_Y�B8A�x���1��!_`���9ê�����2y(;Ӹ|Llj�#IS��/7���F�#̴%�Tx�'&�\	�"�9��W�g�U�-H�y�M��:�nE2��׍��3ؖ`�&TysM�L�����K����b��u��$���qn�2[0:����Z��P�7k-�@F�]���+�z��p�פ��X)��"�L�*%���K���C�� �B��bt�$O�!l�X�SR`���9�w��Q�cҽܞt�H�Q0�r�y>��}�l�ek������_��A����hR�a�`���>�)Q�����I�9D�� �j����K�-#�f���IH9Pe��K�����%�1~^�H����)f?0P�3d�j������`�L�����4E5L�p�'�ĝ�?*�2�Xh4� /b7`)k>|�ݦD��|�ou�+�ŝ����0
Z:c��z������Ƥ��+�R]|g�e�k�l� ��Ȍ�4-~p���㧞{N�X3?��	��,]f���L��v$5A�F�^h�8�����s<�Y�<4��:�$9U<.�,Ze��%}]�<�:,�h�����ٷ��[*���L�)ʫ\�� �Wy/#7�?%�#�{�KUrok������J��{w��#uh�-i�ѧ�H5�'������X���ۍ�>;�Z{�v�D7�����=��Y��4�eg�V���Q���!A��Zz0h�?IH˃�/��AO�f|���+��@�c��l�	!'n+�πȣlQ�������>O�ɟot����=�3��; =>q@��w��f���H	�b���P��{3kU��D��F���a�DV~�1z����uZ���t'�	�\����.�+�#m�����8��e#o��^~V��9���˃-bJG!��=<q��E� B,Z�{A��:X�S��S�?�k��l E����@�t��p�hd'1�O[<;������$'��ׄ˝�^��zց*^@�z��E�s�A�*��R���sGe ��[��kY�᠔,���Kd��f)����w}�3�=I�p�l�ڢ�<�l��ӃZ^!2�%&4��Ґ��V8�o`�>���O�u��r< ���� ��6ό1	��L>v~O8+UE
P%d���D�H�	m��{�w;9��fDd+.q�d�3��9�C�N{�F$$&�6L���7�ک��Q���7j9|�%�c�F�������<���4XZ0+�=!�&�	��[�rd��c~�i��K3]9�^�َ2n^Kd��t�Դ����Dk�v���$H�A��D_�3�|���$�h'��@���s��:�����o^݀h;*�*hPqҀ�x[D�@q_�-��:����}$����Ek�=B�"�Ь���=,U3Hֵ�6(�sTM�d��g��l]�D�X͋�,�J9��Q��q��%�M	I�<�2Ē��ҽz�ʥ#���W�c�-N������G�6k�6��w���5��A�+��?�?�aS@l�	�:�=O7�o?�_����p�L�\�%����{C�Ey��F}��"Z/����N_���#�����{��e��v��r���lvk \�C5�R \�]k̐��L�e��Au���F?�q����gْr�-_���H�!�=΂C���}�����*��[�uiVxݥ5z�_�9�2K�$�-)G�a�䁁UBI�z1@�i�H��Vxc�qR��7�yx�"�+ޓ��Xu�Y�#J}��e�!���w�U'݅p�C�0��C-�~�u��.��j���SX��R ݧ���@2讠��(R$�\ε���#��u6��x Z"?�i8�dvޙ�\�v�I��!��f*�_��ʊ�^�11D�J�sK�� G�*41�P���.�c\���̊�2��c�ɬ �p_��"���F�WA����-v��n�hC5��<�����U���:�~����"���%��ש��죁�l�@g�,n�&l�]ǟt��aj�S� 4)2��UX߿[pAI��XOKR��0��(���@e�
Az�Z9=(KI<�N�!�x����%�`@��uC묕+�߫d�J: ���*á�����">`�t�j?-�3�b�����톪����[����ln�JA�"Oe�#A[�~;��~�}AG�v�[z�Q��^��R`p��:��u��+- ��@Ƴ��H��]�2�Y� ak��|5FK���9�����?)xI.��ŵ�(�]Mx��$~�pGz�����Aoc,Q'q0+!b���哞��,�P��CH�DMz���h^gi�(c�:�ٹro
���a`#����>�)� >�eLՙ�3!������P�H�����h�K����|6j�^�����ZK&y�,C@��7J��+0-;�k�5_&���!T���x�] \Y��l�:y��Ȭ]�g䐧�y	<|��iF�2+�Z��D
�fw.��z�-�J׽9f+�n�mth�[
2�~�����Oen��ϸ��#����K��]��"�]�ş�"G���˝W�H޴)4*S�?�8���S(:�����v�	��)$�bBt�M D�	��Ay�n��h�o�u������!��:d���UܷW��@� wov��$��H�QU,��qOH0�8�.$o�5��<�YT�sX��m)�d�ԿU�hr�G��&FJ`�}EY�f[���cI*����iP�>XY�m���;�#�+��W8r�
�eQ�~�����R-�\]Sr�P�3��w��+o���� �D-Lh�s5Cΐh3�<��U����,��AI��' �"/�,N*�$�pn�+_��b�����Ej=�#�8���?�T�	�S��$��B[3W���kJ`�D�Y884���2�l\�L�a�VR�>��,��va�j�ieY{���Yyؚ��{Nm����_���$B�qr����v	3m;��*�E�5�#Ul��&����"+ʵth���b�q�o�T�X~����eb�T�B����=y{�%����v�,u�nH�1��B�A��Z")'\%E=�<^N�6��7��� H�������χ���!m/���=��_��u���/�z�y��t��L�xF�<`�HC2�������\N�v.g{���+��Rw>�����&�\[�����L!8N���<~�I,,�!2��O|������P�'��l^7k�-���gxF��6˷���B�2ѽ�fg	��WT��lc9�4P�o�$j�� �U��}Mz��{)R��J. F�!�A�0�q������BC����84���Ko�9$�⧱��|c��?jK�3~к�a���W7WR:�ס�ƃWS8��0���sz�ϙ����PR/�u܊��]$���O���}u��0�F� ý���)�6���q�����#N�������(1M�Y�Ӌ��7��+�xp;�4�%�^��s�k��+��GnY] �z��SFY7F�z��.T��1ws}�p�Ű3s�/ ��W-���Wj#�MXZR/�V�=����~��bp��*v�0"7��ٱ��b����N1׿7y;�T�q��Tw�vU�>jL�	�$ϊ�C��$	|��^4�oUR�	��7�S5�r�8w�.�Ӆ�Q�߱��0�gd�D�R��{�N���_O2�� E
k�ھ>��j��*1ԑ��2�+Z)����V�}�݅'/���y����qu_��꞊S��Ћ4���-��ka���ΝЭ1�^�9X��������?�ł ����+�f'���'�8��L������FP�n����((p�Ԕ�Q���dO�cG��6D�Z閻v♿�3��N�%&i�XW�/avVik��P�χc��8��Bfh!���buP�XCw�7�-��"<��&��U�=5=4VcC>�\��{5X�tS5'T��N �X-EFy��[�XBTjխ���/l���� ���c�
:ǿ�-� �'&����# �Wȸv���e�r�t*�=-Q�@�m�+��?� =)��������n��
�2L~if�W\��m�$����D�$�]�p�&D1d4�_�K!�����G�ݴ�C>�#w���$�F����������X/�R��P���M�Oݏ(]ߤ�EZ�g�����]?)ȍ���������re D��SAG�-L�W�Y��Ȫ<������8�*�J���Z��L��F$��lj�)A�&�Ԣ��f������p�o��t��:iͰd��䵌^D����_u��������f
l�T]"�Y?�G�d�>s��qWİOK�`p3�{v���
��hgJϫV�����{�Z�����y� �BL�,m��f��;3������a�I�0�>�7t��Y
d�T��;0��op��sL�Й�SR�?2,Z�P�.H���M�����|Q��֮�&P�Q����9Y;mc�����-R������C���ѧg��m��aRP�ڄg��.�6�����
0�'��հ}x���I�ě e�"�BKs0��V����ﲠ�Y�0gx�ħ8��wv��1��~�q�y`�8K^X�)H�2y� z����(+(�F�&�1�(�'����x�%��i�Wi
H�\�'*��߱�����@�M^���G�"������i)�1�#p8ş�Ž#F �k���Kg-u}}�n@^�"�k��4��w̶��g��s�t<����l�N�"l��P���Y���)�JF����9n$}���LG�hM5�eR��<V10�D��,(�IS��U��.�~LJ�x]8FQQ	lL��t�t��5-�2��fް�f�	$�Ģ�g�:�o�Ktnt"`��̹cη��	�1�7��N4)���:��U�(�JC�kn뷙�d_'��
ŋ��~#�CgA
Qo'�ZVu��7X֕a
r<��@Z�:@�R�.GL�a��ar�>'�j�Р������Ӱ>^ �20��=p�%i��z?�7/�#m�xB�$$mߖ������LE��u&��jG��/�X�}�5/�3�D-�K�z(d�q�X����9O�h��f�r>�SB����ؑCG������tĸB��m�tn�$[N[߸x�Eס:5���n�[SJ�6�3DWn JAGUa?���2$��[�~��	�[�fA���}]�EC�F!��)M����d�<t�v�|��Ȇ�tO��1���ݻ[��(4nyUHN]�4i����#Җ[)�q�x�1D�ۡwij��*��;�&���i���B/ft�����;=Va��u�4�X}��
^Ga�Vm�G�\&��=�(>�S��Z��v�k8�e�C�>e�ȱݪ5���`��y�B�w���>?z�H_�CzӦ=�Y'/�	����/�p�F����e�n'�>��v�k�1�Z|��	�3�#�Ӣ��/��Po�d�W���]���x1��fq�5�[4�B>^�4��u�0��{թ�M�8�F�+Eͽm�4%{A�:ֻHv	GV������/Q!_/J�*�Î�K�#�=v>ғ�H� ��kX�����q9r8���"Oõf?)�q����5/�1b�o+��ea،�U�������7Q׮`w���X@EDt׹�'+�?�xE���]C�ДY'��9��,<���N�8���w��9�����SK�Cr��p�)9~+16N-��7)�)7,yt!��h^K�uncU<���a��ϴ��1t%���:�C\<�6��|�� U�@��kg�������,����x|�3�`|�7y����L�jL&ȐP�c��['��rFcn�
*��g���zq�7��OL�,O9�~r1��OM�Fw�F���zz����K(j^��'��N���|P���ÔyH��Fa���nR[����\8��ۢ�Û��Q��Ԅq깍����&��1x�w��s�Te<��WZ
-� X:�������'v!>{^n<��hY�DVƼ��-�Kdf6�=*�?�s�_��J�T�ꮴ��7��Z���%]^����q�2ҩ�N��>d2Ԕ�T�o��E�9̄�Qy��ʪ>��^0j� Z�򳲽��+nyl|����#�/a%ǘ�����XM ?l��A�]��|��T2Wj��*$e�k$��p,|�ye4�Z�mS�a���`fL��E�&O5�P���-.�wL� �h�f<�u���DON�X�{?���|5�� ���^}0��6�f��^Ϥ�����3���[�[�%�v�X	�ZM���D�$PD
�A�]��U���;��`��H!L�~ƾ�u�hi&�y�B�8��m��IOZS���L�KN�Ý�o���/UF�✮�����|L�c��72xx��G�|��5�NBo����*h����b��I�J��WN��V���t����$X�MY�x.h:G����u�:��"��R�Z�_yD��#�P��8IC/*܇N��Z�F���,7W��@'*��S<鞐� �Zpe���_�
��X��:3B�Dg~�by򆚤��9���<�l�R��6�K}7�	%(� ��w!����(��>�bO$����=��++�?��q�J��D'�d�:�n��;]#��"��pn��uv�,{`��U;o�A���Hg��՛P�ӹ�y8��}%"$=|�/���Hʄ,���.���a"��c��Wb�0�LM�ωv� ���*��L7�0���y�7�w�l����8��{����]�x�LլW�&��"��h���/eX��^�.�� �j��'n���R�y�ۖ׺�"�7�KEݲ�P���Σ%Xw�-a8��`�Yg�@����&�(b��d�v��m��My�~�C0�h��j�3^�Azo��K9�{q�����F���$�Ũ�Q�������!�!�S���"s��~;z��M���O����҉s4u�Z��t��͞�c�k���Qel�,��ެy����4>�b�3
HB�˺R(0I�X�;��
�Jsc�^>e�����T�@��}�/&ϧ���X7�򚌨�������a����Ebq��*w`��%U�˥;����J�%�VUgzY�N�� ���\��ߖq���MfRa�D��a`��:���f������^�SP�d��#���+���q�td��!�!�{��s:�t�%�����>ݷz�p��:�uf�i��o��<�1I��f�*���O���0~L:�e\<��?}���ۯٝ:7,�M��1ɝw�iq�9,���\�/�|�y�{H���^���X��'�	�#���w�1�E�6M�e�g����TF�%K�m#8��D��y(��}8�EI���y]���S��4����b��`^�-�-k(|����J���r#+[���*�Z�D�dg�C
����ĹU7�J^nȮ�h����#�9q��q�7�+l�K7��`�~��]s�;�f��>��T<��T��s�)�5�Y{�̻\;HB���y��6+`u��謬�a�m+�.���RF�d��3�N-���-���;�m�WC�V��7��ޝk����K�n��I��#��_��T�.���5*'��t�,0j�=zɈ�܎˕ϒ��{3��&�Y�2ά�_Z蟑�n����<��b$q���^嫡���p����jJ�M�T,����
k
D�ւ&���j��l�Ɓo� 4�8�X�n��;���+s��q�HY����/���<�;,���N��e���lQ�%).������͑�ջ�S�A���>T�w��O�~�wަ��|Xq�LP[�j�r�'�Z7�$�&E�wj��R��OJ{o+�h2w���p��Gs-�t�@��̒SF��|�Y��Iq8WB:���$�0S���T��~*�[o����{�E�juE� Z�m��p�J�	�{\\�1��^��6�f�p�$���<�6I�'/xrs���.�d��4y����-V�a�Iٗ*D���~; ����CV p�o6�>�	l�8;��&>౷�8-b����l(�qq��'W�3�j�L':�s0�����I/e�`O�2��H�"���my��`��DK����?A>jg����}Y�,��X�;���ȏ�/�e���s�a�ka��r�<_7GK1\=�[O����nl���$�e�y�̌+\���LU�?]�}f´�~�Ұ��=`���R�[������O�Ɠ�n���z��J�v�hD0�����{��`Y�w����i�����I�^dK��&�k�y4凁ӡ�8i�?G*4DO?5CJ�o�
�t~Vjc�������G�4r�\�0/�;I����J3>������<K-�$`�x9S�"���Y| ~�4.����I��`qf�[�,B�Q�w���f��'�NΥv�σ2E͋�l=�X�H0jo-��	`�N�f[��憃A�Y��9��xml�<�wLx*󾴕�׫!����݀�qHcFVI!��iґ��h ٛa�`�?��� {z>)�{C�-�w�d��yD�����/���7���ۮi�^�_K��bd��Y�޺�����۠uu��o��O�"�X0�ܠ���*���5b�j���O <Q�x��9���x�q�Rr ��D�X����˖��rv�d&�4\O;B�]:�^�c��1�%��	"x\P%��ī����]ʊ�j7��JQɆ7~��~�º���.&ܭ.��]�r�S�A�*@�I�%�ċ�b,-d:��Mo��9�;�44�ɲb�x* �3YRV*��q�->h|3�M��hJ�l"܆��8L���!�x��W����K��i���y����+�XjAY^��x��8�4��bU���M�	aw���:�6��u���,Lb�E��۵x����Q﫛x�`�l���1���b��AP��0[~yX��;+_ۭ�%�-<Е��)M�r�^��G� k[��+�1B����ė��,x`�0���^���$�����K#� |� �MMz�j.U�j�!��Z�`�ˏ��9X`��9}Z[�, �(�h���#r�q�a~��&h� �}3{
���"�@f)��ϣ`SRh�"W���i)`�u���_[�c����,��R��/{@h&��d�$������JQ������FsI�T��0,X��f�"�K|�(% �l8���rCh��a,M+xK�;Ay� �xQ=h\k�c�x!*����ˤni���{�x^F}P	%g�7�(X��}I=P��,�|4�f��KEe3`���%�W"w��O�VaM�3��#`9d�8��?�Nb��i���w��R��"eû/����%�H���g�+��%�t��
���	�H =�l�|M�77�E��&��y9�jǉ+(�yT\-Hmר��u^C�����?��[v���V�8,�D7�D��qG����͖'�K:��ܞq�q�SFr���a���"+ �1_#[��E�YFc��2`*��Kx�.1�*�h����\�Sv�`��Vʂ���� 1_�z�����x���{�����Kp$��ҳ������ܷ´`����UY���7wW H��J]7:����Vܷ�90.s��7��'ΓO�O���h�Y2�����m�e7��4x�#�p�3>JOw~�?�½+@M,�^ �#�#������l�kM
��0��q���bm)�m��1;�?��3�.l2�Xt^�����ˎ��������k�S�N��m��dټ����rk��T���_٘(g�V�c�Z5�u|��L)h�8j6mߚZc���T�>�_��7+q���]�: h ��@|2��}�<��1k��O������s��#��7��uV��=��J��vE= ��C��L>n[�÷��_;�f�v�T�qQ%C���KNp���"��[��@WG<�!tY��"%,��d]-�����ټ�䲇��yU�?�X�SM�K���͞�/�ƮKB��R��g�֦��5���_r�J��C8�,�o��R��z~h8I���dS9�@=Љ���H�=���f`)#���S��ZK��lA@a���!��v^�PR7���Rw�{�T��r���{�)���X,����R���̺)L�.���͐��
�eQ3G��s��h^8퍧V
��W�RX˴�)�<�q����� ��ل��h_uDޤ � �9�#x�h��v�v&�d�����M�R�����2�7a�$B�[�jaS�_M�����dQ�W�O��.�5Q��Ee`k�ኧT����q.O��1\p+�%����%����@�1)l�0�_�t��K6yh��sJ�JMOHOYv�K�B'F��%7�-��`��X�p���'����c��b.�[_�ᯔ�!xiǛJ��d���5y\��շ��$��"��v�MnX���ۻ���nh��`� 4^� ��o�3����ۼ�ߺ��5�^�,��11t~��L��t22�6ļ=�����Q��lF�h۶�g%�?�j���+7���9#7 P��jU�db{*�;���9�K��Z(�B���J%��@u�zt��l��$��x��Amm<��!e��=��/��x�X�`���'v���Y̚V[�ԩ�Gr�(\���U�"3?����G"�ǿ���?֝dےȷJ�Z鍠E�{�Sb����lt+���,�Y;�f��j��Y3xVH?�z�K?�p��n��{�*�f-?�C��f���M���e��i�ě�ib����X�������h���ozq���i�X�w�\N}�7�uX뭎������Ƽ6��%�HYW��&��j#��f%�el<[����KKp��#J~w��B��,!��ỏ2�9�S�"�;���O��d�[��c$v��ض����?�d�j�C��y���}�q�w���o�	̊�午��3y��EC�HC����k�vk�l��An�uN��f�h��į�r�	D:���(��To�1��,@z��,�b���Y�ݻ{�H��s�*"zR�>����U�2�3�ȩ�W.�oa�&2'���퇙(�a�H�F{���7x�sZ�1L�B�{��r�'�H~c�]�.	,~���3�Ɗ����<���3��!���P���W�Z���#�Rc����8v�N�}�`�n'�eĉ����>���-7��>�"�]�@����,s�cf�c�!Ε��(K�b���.C2�c>�9h[H� Q��r�%�}��!a|d7�hz�5̍��ٸJ9_�GƆ�qg�����N�j�O�M>���#�j�C��6��X�X�ǆ1>�_Hl�V3�k+�f�ՌIO
$�+��c$$E�^�g��i�`,��	���9 >�}�Sݫ��Nk�e�68��/Ki$�5���WgS�O�cIP�Mk�=�����ҐayZ�0�&�b�}\%��#�,��'Iս�@�ӄGr����I=����L��c�@2�>?�v�� �Y�v�����HN�����9T�l�uA���Ҽ�> ��޹pe;7Ҩs�'��H/�Y�~v�	M���בJ�&g]|�A#(0@�P��S�`��:[v"��ƅ)�b~A��0��^�,�A.ڬ��Q	��j��E$�o?�S�3�=6i�����9�ҷ�{�0��(��C��Y)I�����Z�u�T�7C�A�u4�L(�;�!2}>�&�+LU�+�pYuvG�y�I� !>������,���iԮ�CT��o��P|4�O%��X(�s�`�}S���x�;s䖦^'�w��zW�������Ƭt�wP���v�A��a�y�n�Ϭ���ȑ�f�!���UBqY(���Dj�Q�p6%Iu��易���"��1�g_h�b�_Mv�j�P��~�������L�=iO��EG;mG����(13��h,G?g�@�p���c��آ����b�p��
 ��w�Kx�>i��`��K7m��Bq	/���-`�����Q=��	��<����c����+VhL��$F�/��9?I��OM���ۭb���X�Jc���;��-`q�X��JMI+�F��^(�6{��7<�u���!e�5���x2�.�i���d�{o�/�A[�Tb0�%���\J����fD[C�\	n�i�c�F��)NM$O#���PEV	�$�-1%=��U�c?z�~I���cת7���F~+���=$T�9��\Γ������RZ��Y�(���]O�As�j���Bb�<|%���ҁUɽb������@$mE��w�Ge�Y/���$�q_�:��D�u���̊��_6F�r�L���s����2v��G�^�D�ҝ�Oݙr�kZ�U?X;fy�~�O�*%�әs]��p���A-am� dxA]*t-�q��M��i}ދ!/��i�:�)�Y �8G����z��ӡp���w7��^���s$t�|�Myr54礽Gb�L��Ĕ��N%����n��[))�2P�Ҩ?ZH��W�qx���S���b y���<��<u�'Ql���!�ɽXq��m}NE�Xݑ���h�:v?�?��Һ>�����0�=�/�P���E1w�:Yn�
�!0O���}������-�8��~�	d�z���E��wd�
�A"�("sL,�>(k����c�@x1@?ug�oѼ�K�3�^�3g2BZ��A�`+c�6� 3b�}�)���P��h$$x�Ȯ{G�����V�[m�N�n�eT�{n�^X���"�<'�e�5��?Y)��=oE�d�uY�y�ࣕ_��(��J18"�X�~`����L���}4Ȇ���aDVcw�
����S���?&E��4�slT��B��d/�;!���-9�Ks��B��X�,(ʑ`�J>�W<���������ut񽗏7	��}����2bO�?�b���>�e�����pay�=�?y(Ml�lZz��0ʽKY<�!1�F�}+ثa�h�d'��Ŕ�z�mWi �+�>��{�F�5��X���1K�t��WM���C?B�K��"����GD�o�m`KO
��O���5����^�W�O�#��m;N㛲������*e���h��$�q��u	.:��(�_�a&엝�95�vP��e�P]�$�O��6�Tg�����ffYj,�Jؚ̓E���F<ՅŐ���_��ؚ�OYzĻZp�D��mJ��̮O�1GѺG
��pcB��0�m��o����~�i\D�l��k�s����r=�n՜D��,�b&*(���>=���v ]�8䉁�P@6�:�`9߶z��^pk@�t�l�0k�k��hx��� �f��.���g�N�����U�Z�Ժ��ྞR[hoZ����ʁv�zDmx�챮\&�kW��&S�]�k�N0�_���r���@d!Aޅf
�A�m?'j7�I�r5�MI�J}1��������4��	�ԳͭA���ꭴ%x��yDA@���%R}�&VZ_z)H%"@��O��# x����´´l�TC!T˗8!	�;&ź˾���v/�p���{޳���������	��s��dh*t��a�^�3��8ڷ��T̄dj�ѩj�V�uPR~=���f�L�?zU���Κ�*J����)4�#|�p7�Ze85�r.�曲b>����q�N��:��ƻGh�\q*$���<����my�SI��2�!p��F�h���(�95FA4Q!k�ވ5�I�)�Y��k��~��7�A��I����U�A�Y��c�)�]���?Lg�E��]�;I���6�@!��[e�DpaQ3|?�ځ��)o���ޓ�n<N��2���WJ�H���؎��ay�L ����D�i�u|Ay�y4@��z���>Ȥ��x;���:s�_ -�_8O��ܞy�0_����n����,������Nq�
���yk`�y <";��AC�K[�g�Z���A���y�'a:�Dmxs'zDf�g�k-�m&y�Jl�~��eG�q�.gU!���UfA��K�fP�"�
{UCm�ҩ��� 6��FV�Ĳ}�
l9ł�B�������b���mʫu�A�ϑ,@�����j�	^�p_3RYk����˻h�y���s٘�7�{!��&;)y��ТQ���@�8��5�[S��`��҉�U ���?���&xgJt�4�c�#f�o��Ł�< :8j�T�a�&�}�R� }�������pȼ�6]���d��v�X�J����M���b�T�xB�d��ݓ��[?x�,�Ԉ
��� �j�2c��/z`��C� �T����Ht��s��HL�gab�������a���������J�����Ʃ��C2h2
�p����J��UQ��_�v��������%Ӎ����^,�)�>ܐ%�\����H��MR7�����Bf���$������(�_$Mv�W������-1l�����A������s�%	Y�o�>2Ue�І!����(�Mu�Jeo���� ��m��q���%4��L-H4)�1��f��h[ �8�P��<�sַ9w�p��B
V0 ���L��;�QZL������E�ɯ�k�M�3p&Ѷu�O.1,����^�R����\�cךs�3z�-��Xp������5i�
�̔�<\�ȗ� x��&�=�d��}�`3Z�v�����uX��s����fN�T����t�/M�Tm�53�*@�@׎��K���F��ث��������.iq�,Z����	<�
V�,<�������'�͑V�1�d�0�v��<�,3-��C;�V��LPw���?PualcP�2����7x�/��,��y�6�qn�k(|v�Z�A<�Y�I���X���lT�x�?�ф��*�X�:?Ċp,�2�4@G�[���ƥ(��-:���%�	xj��?�?�Qr�B�Y!���*-�:e��D<��Fd��Nh_�*����ݜgo���x*[7��UZ�/$l���|�]�+���<j'8��)܅K�y����>xpܥ���	�hm��Q'-[�יGXRA�̐8䂦�'ڄ=bWk b9�"���Ec���Ic���%p��vub=/���-���s�l�@�l
���q�����'�~�� �B@:��ڀ M^���$r�1K�C�����K��"{���+2�L5�E�X�?��}���62���F�·�WjB	����D��m�4.=�5u���/rƽu�ࡂ(����F����<��'��r���"��w�]�H4 ���)\���L��ґ��k�_�2��\�[�=g4�>���w6�?@�Ӄz��)�dI�Ft�N{$��8u��
H��nl�+�~*6n8ۓ�L��_�zn�X)8����g���������W�����H���]	�z�b��<]�$����UD�% ޙn�{���~����f�o<;��V��P�
����uX~����og��PI*�y7�_��O�Ö��¢x�dО���Qcf�װX��;˝�^=�	_ ��Av$v?{:���_9�|��*�`@7�����.Y*����.qJН��]	�h�Xӽ&��gF���ok� �s���}\�~z����_�B�DӺ��4Ն���L��U����G��Yc,~�J������0�6/GB������yzP@���q�����h���Z���|Q��r���`[��%�ë�|,ݐGG���&6��'Cl>5+�^v�;����:`b����E�8WY��{�X �5R�}t�~v����1Du93iÕ�ψ�JX�r����4�Y�'	 ot����-�����=x�+��P��e0ۄ0�=�/�͈��C�H���'�ؔw}x�S�J�c�:�,��H*�rԌ�]A��~|�?�/��Y�^��0:�J�g���G���DӘ�.﹝S����ϪL����/���h�����F.\�HT���2�kx`W�GJ1�gl.��GW���>8�5�H>�7�6��u�;C�c����������	�%mE���ˇ��̷�ӊ��R$���C��C��DŔ�YcJo$�p^�%R�u����Fӎ�=#[B!�"��c�]��O�[6���BK��k��>S��&m���L�`3�$���=冷��� ��n;�;��A��l�)]=_y-B�?���8�����Z�u*w�m`u��c^w�{/�ʸ��&���s��}T�P�RF?B��w��p@"��e��<���&�Sj�T_φJ\{��w�^R���΋o��Ռ�w�J႙�n��ay�lk3�K�៦Z��Dx�b��v�4��ϗ���80#K���	4���6��Ug@�A�RY�{�d|��Gvg��i�I��xX����b9W�0�5��WR�W,�i%I�I�T�V�tZd�c����ph�'=��;�C���[>�7�8�I?t%�O��Uχ�xh����ܧpV:92A�2I�b?�V�|��wY4ilA�=2%s�����䠣�Зѥ����Q�A.�<�ĩ��8'�C��d��q�FXQ8di:��/����>	�-�ߗ�#���!�X�\v�UW��������S'V&g���dT�5�ލ�f�3/����+�h2ޘMzY�Y�ϊ����$7ݩ�j�q�����������0�,qj_V�b�L-}fѤ���+�Ĝ�@��.��)T(aJ�$=�D��@� ��37�̕�`+|�q*�����6�=�瓺VqY�5��!
&=��+=R�r�W�j��AL�H�GP�V"X)i�����W�[o|����_ZC&ZU�4�顦��e����$xc �)�A擄�z%P��w�랞��Z0N��c{s�W2�_8^'��d�+x�	�zx�Y��X�Vrq��i�88j�YR�+$la`:$1�P�w)�,go�5�IPHV�esVV�C�[]��Lr6����_ �c�!UVT)ҋo���uZt�5��੕-�ќſX�w�5�۳�j�m�CTA��(؟ZMǒOi?|^7���6І
O�ۤݭ����=��H���\&���q`�9���;d�ԡ��1(�T�<�7c����A���9[����k:At讏��陥�*�.ͅ!o	�6�O9���M|��WM3�\N^b �C<�GC�9ੜ�����cm�ѕh��I��_{�~Y��� �/���@��ЍI�0��e;��ƍZ��w+��!�FȔ� pԐ`�0��+��N����q�~���>f�sqo��빯�j��oyY�����}���������_��,��:w�;Q�=�������
[�T�1u�>�xm�^!����ztD��Dp08����%8��)�������I.g��x.N2�tm<�Dt�Q�p�+@��lw�ڵ�9�)	��J���h�ƙ���-����(o0�6p�Ǐ�٭��,|��G��l��WE=�t�z8�E�<n%�Ǳ�s��(aTH�ޯ���e��_���6�t23���>���FO0����I.�0X4��0���fbh-�`b��9�4��v���9 �g�5�?&��mRmy|@#{.	n��Ne�*��L@�H���\�w�����pq��/�셎Ò��ê��"�0XH�a��	�5��)�p�[�0�'+��{�_ygǉZu�KJlH^F�������3G��XM��l�;����ŀ����[����栞AXtȉ�M�6"8-�#c㫮���x�a {���A�uOZltS��]	
yH�����1��ݽ ]��y���9Cߛq�!m:kƝ�[S��H�G�!�����7�g}Mtg�}�͔����P���T�	��{\d��vj`�L�h��X�]�6ķۊ���k�t/.%���sM�v���G.��8d�R�qKn�(�A��@7 ����G�'��{���Z�.���	� ��o�P�fͪ��*��g��=��$%��C�;R�0��F���I=���hU�ӷ�\�m���� 	����&�!���Ղx�d
+�r~���E��㶤�o��o垝X}-7O��5l����@X�֐�z?�g��˖H㙱�)��:ʛ�__<�0��t�v����!����m��;ŭO`K.�'�z�BG�ϣ��U�fqY̪�+b�ۘ��:�w+�8_��`�Yw��ut	��'1�x"��mL!��"ɒ+0�&_j2�R�n.P���}(�NL�d�L�o�<��J�p/�Kuz��Xa=z�(M�{�_�k���bWle�� �ك�l�W��ϺӦM��������������r�Q	��pm�\m�G���*��
��wNX�@~��݋�!I]2[��|Uq�.�NK�<3i'�|G�Y�h��y�u�YH�LL�٨Nb�"�X�3�p �5%�X�r��Ḧ�H�\�e�+Rʭ������-�d#�b�/�Bę�Q�H�g��);~qnyy&u��;�`W`k��L��X��,}v�u3a��9���xx�?�
"R�d�����9s��6���:a�Հ�F����G���|Ǽu�b*Zy�r �59�HR1fd���A7����+�+*�Y 硶A*�h��`&�a^�'��\��n!Q�.xH�n:�M׮g�pu�c
�_���\�o�q\��%��M�[���{~S	�uz�0Լ��@d�+m^�X3	�؀�p�"� ]�,^�\��yY���P�;�v��7m�!���
7�A9�dm�Q��h�h5a�;��kϕ�����c�e+/asv�j������j���,9HV"��d����z&p��U��Qv1q��7q���![�v��K$�VR���s�+�V���90��kX��۽�:ߴ�1W=�9���!�^�O�4����ȴ�p����	GD�P����6���<�F�(:h	s�����۩0�� }��D�`�N
�5����&�?K7�]�D�I�����5���H#C���W��δ=g=��9�hy�3O�	��r��%M�e��*w&]��e�#6��z#D����7g̠����t��8[�2m�Yٍ�m�ֺ&ѧ˦��w�k�
{����P������2�d�f�#���n��V`�n4y�K�S���1�?O�l�2g�44LC���-Va�]E�Q8��񜤷0�ҨC�;�O�_��⣡�6�;9ad��u�z�v���U����c���L��t":�ŇJ ;�m�Q��%e�\��U6N�:�!ێ䵧�.;A�U��oc���v $#������=�(�cVOƟp%rTsy��bԙ���������W��B����Wќ]��^�Nk�a�&��>�(�D�
j�����6I丌8P�S�&�Ey��
sy鑀�������<V�UK�؜�<	'ڳ�p����*k6��N�HO�}$���7�X$~��]�5s��E���)e��g�%U������;�>�t��j�z�N�	�!K�zs�G��.�qK<9��1��4�ρ��<3��V#��@��{�VmS��:i��7Z�4�{�d : ys^#x������a�֚���x�*+�9��bo�:F�V�e&<�a���TM$�o�
%]5�u���'I�t�<�D�c������^�rE�s�KM�B��w����ǒ4��F�"6?֘�t�3
�Z1KR�cn�C2�Ţ�H���bI�#@��Ǻ�ȯL�l��y1)��-R(�8\G*-�Yå-UF���Y���n:�q��X����?!� �b��50�>��v�62�'/!}/vI�i̊YǕ]�V�I�[.9�����(l	��|y2j��AU�D<��|bw�3�a�Aá$��Zs`���nX$�ľ��n�jT���/U}Y;#��*�{*�o��$/�+{��ڻkˤ�o�}�,)������K��m��Ѻ��̅��]-uX丮`��5"��K�{x%�5G�	����e ��L�����	����U��)���_R+(�<��\�	si���駎=|~�v����A���3qx�t���P����x,~ �aU�r���a�-u����:_N��W���'R�5@s:F���r�*��4J������f����!|�����t�(T�����'>ۄC>�KP*�����1�����H�H�ԡ����Tt4��k��0���SK��
V�[���犙�N�C/Zu�9��^�J"�Ra��A���Nc��'8۝#�~�G����R���,�r���L	��u+N''��8<��4�ܟl�;�G�*����Zi�o�k�ߒb-xZ�Qp Vn��}+��$�t�c��������ۊ���4fg��m����������-
�Ф(�)@&�Bu+n�|�j�(���S
���P���[`\Jmc�5�6�P�}`�/ I����,�էp-U�H2Ow<�v�����ʣ3X���k�D���`�g��[���@�m�q�|}����Jp�a ��YN���;�Gp��w��H�����+���7��o~��c)9���16��BŎ���u GVw��5�����]���j�h[����K��B���ib�ёH��wVF{�Q B)M���M��'����ǝ��7#m<��7���Z���_=��:֘=�R�`+�����r���������|	]�@���^�r���rj~�-t4g�D#a���h�`9k�Λ��(}$�%��'���q	 �_����αj/)-"��yܒ/l7�6�f�΄H�§����-P�ۀ�{/Ƽ�_���'�w}��� �ٰ^
>kt~pS��R0�b��پ�mb�r��wo�U-^�vb������A���cN9 tֱ����.0���\�!}r�����H����~�\�M�����45�p[�~#lgv�DiQ71�<3�SBZ�{ȯMKW�J��@³�&�m�3q�U�\����a\���r�`}u)��OQM�;�\�I^r�8�T���F/���#�[���@��([�����U3�fW�X�bs�bX�g���q��Z|����g�R�>�ZZ�S�"r��}��耰BI+[��7��T��ie=�<ZaP�_��M�)�9��5\�CG��xbþb� ��x ����j�I0u�5�)M�yM�tg_�����Y����U*�1��:�)v��#V7o���ۿ�Y��*}��T�*�{]��n߈�A��Ba�D�Z��N���S�M��gA�\���!���0���j�Dk�����ƅm���;/Z,y\��2Q+t��ˬ���c�2qc��;��))��T�Z۝SIdf�X��0��4��Ƃ�FB��c�}7��8�6�l�@��yg~B��WF��c275lt�q��z͛l����Y��|Ojb��b�U��AB��?�o�>�>t�ɀ2J������d|�ٸ�(��o����L9:�먣f��Ƀ*��+)&�����9&q,��t,�\ʏ3�i}2�s+���S!W	��ձ�}[��>tD�zG����1a	bm��h�'��pwGّa3��<ly
�+aN4*t��g��Q�[Q�Y.:�Ŵ�?�%�+�U��oq���I�aIд�^�A����i�r"�C��m҆ ��"�1a��G7�W��`*(�Q5?�����0�7��m����}��,~��2���Fo~:�bBBp	u�5۞�P&Z�:_+���ʛL+���m!8&:���Q�����JY���zU���eda�q���B-����0�Xё-�ϊ�4{1�3��͆Y�s��xp���;���ͷ�RZ��$����NS�&�Hܔ�1|� �4C0����}c��C�����zm�������r���<�����X���I�AN�?���Y4�2���Pv�8C��B�SE�u���8$�Gޗ�K��?�����z��}?<w�W����ZT�*6A,�v��p����s�#�Y��;����SJ����={�a�9ab>,���IͼN�> �"bg-8�̎.�$��jW�_\�?���՜��`Q�<7�Ak=��=a%;��b����C|�����g����T�	����}��ov��*�w��ٖ�^�L�ҿQC84,QzI���۳V���ஈ�]{�?Q�f\<�0LC5�����)t��2Ά��H�8�{�f^��#��w�
�摎�����x�63����^ͻ��8!�s���ʲRi��fs��σ�@ ��Q"1H��e�7���g�p�ѿ �� .'+{!�7�=���H�\��v�?/�h��0UH[�^���k�"�cJl�M���Б89|6�;pH���ƿR�ȣmxx�����7�`��9���	�g���Ӧ��L9������Jݢt�FM�#����\��w0�������@cf�Z�aV4e�.�H��Ú�k+�6�I4ѨM�cl�x�1lb7�M cB���q$Ɍ����E���K��,S���GT�w��<B�S�JD/($�Ty�\��ũt�i��5�#�A�7i΍�g�{�߁\��8���'(ۉ��o�Gt�'����ψ�V?�)��g�N�v����4UU���@����V��-��.�$i����]��	�<�2Uc,�����7�sG�y4�����A2�F$���L+������'[���2�H��Ƞ���I����8gf��#��KX��)+���<!-0{������`�UUޱ��#���	�%����
��a@7#���r똢"^T��
�㝳 ����|��;1~u�y� =�KS�چE�CS2�+8�p�����^������J�zJ��V�mZ�!ZR�u��	n��z��ȝ!�=ă�6�:�������Z���� c���nF����I�<_D�#��W��"����Y�a*�����	��[�����I�����!L���m�c�'�*��Ye8����?����`:�a`��t*Ȯf��Y��c_"����7��+*���pPWuc$�".��l�	悺=-)��rey�@B^F:��/0<z�T:�v����fS�x��?
�{�o�F�_#W�_�4ˬ�p�(�Nn{��e�x�cB����Q����l�c�	�������
@i����`�B3'ttf�����n����1�O��!	�Oq��^�Wj[���6����/�B�f�'�ê<"���������@o��</���R��W
�ι�2�`���hUg��^g�_/��i��hy���ⷽc,J�ֻQ���O���� �}���Q��\�3�J}����m��Ԓ;œP�G%���d�O�bZ��(���N+Ҁ�a�$�S����	&���R2j���,�����h�<Z�װ��EE�^c�΃����(�^� #�<��C��6b�chO��_0}k79Tq���8c�z��� �A��&5��d���c���Ps��U��D� YX��P_Q��%��7��f�'�R�	ˬ��7�/�s�kz�����	�ᄼz���j-?���N��y�)�{Yj����w)E�Y�AM�GM䴤Dy3�ɗ���ӟ�tmo��jevȃtӄ_��3�1w�s1P *W>2~�"�Q&�֟/j����·�"{��A%0B�����DKǺ�l�Ziʆ�l���ʴ�LP���� S.a%�����ڮo�\�K =�|4�&1r�'���$|���� \h�3�s%B����#���x�+byj�rBZ���0gF��}Q��9���V ,�,P*��X?�q|�E��=M��p�9����eW������*CSO}pn3��ӌ���ͳד�|��.^�x
��,�ף��.�������VTK8\f�)��e�������P�� B�K���A��
J%čs���RC�9���_�Hvn�b�(��)g��U�e�w%��%o߃�Nw��-W�Ψ�G�ޜ.�=;R;a6A��&̏͐
�p���ɥ[�0������Pk�
v0ٹ�z.c�� vV 9`\mZ6�oN1V@�(�ޖ���}�ޭo���ވ��G��0��19��p?)���9�~-�i�GG�?底��K!V��-�,Tu�G�U8|}Ml,�s�����9����pK�F0t�
��pn9�G݌J�C�`)�a��8����qUv6�9��.�Io5�D���<��5I޵m�����t1P����?n��&�X�&��f�x� ��,S�ȵr_.�RVt''v:�������be#���ېb�@�ת�gWڈ�t�& h2���o��OC�uhu	ܼ@E��)�{^�ezɕ�:�k�JjWTtѲ�?�q��h&��<������ݓ_]�7ȶ�vS�$�|U�x� ��ߥ�yz2~�����tWlp9�Y�~�1^�4��C�})������i��� ��%@5�����HG�(Cn� �N��)�T''Ww蛓�����7yg�&��	e�v�f$Wmی��T�Z����Ϩ`�E���AO1g,�@`���ީ�r+(i�]��)#X�n����z}�P��{?�[REx�GcF��{2���n��},r��x|�8�5�i>�\E����Y�>&�������b	����P����s-FS���x��|�Kfc\��ы� D1cF*�as��4�F�����rv%m����\&���3���r�M*/���������w�¥>��G����)FC�_����,��f�#lXX��& �"�jϾu�q��L���rB������z�>��%�.��pTz}�4�S��\M�&ep�l(�FC^�����c�fH"��>l`����Fq�$4�ƺ#�����[ dޫgep��c.��G��y�
�����m��5�����B�������'L��]R��;N&�EQ�c��C�;���<G�VUJۂ)����gG���#~ӌE�'�����p^x'.fz��39^?��RaL��
h��Fe���4~E���VG.�N�\�V-�i%�R�IX��>E��/�.�G����0��:��͢d���>6TV���tS��i�d���7���z������6����mߑ�4T���x�����د���hʗ
5��]��#��E�@A۴��/=�|�tu�ś����7'�!4��WG;/b��;?3���A}.ȩ"rBoΊr���_�G�hZ� %9S��fM���y/ϗ��bOD�[$���_	�X���BV�j��v��1�KI�����?}�xT؅�rȂ��~|�v'Xx������n�2
,9��aX�g����j�
4��Mq���)��t���Ij��v��W�XA]�(�\	z���D$�����&w�2:�.qL����m>V��*Sg�	�aW"�JG[��9�4>MJta��Z�Iݟ% ]�5�X�ʟp_�b�ە��?��/N��4qc���X���JE�W�3n׺D6� 6О����([�:�H���z�=',r�J��.�31���'n�-{��"@ 	"���B�5n}��ڰ���O82���ϋ]���6����('��Ǩ�#I �3�SĦ��[�U��UoL̽�����p�H+���GO��m�:-��w(3K�X���IpN^��Yy���&���_�V}�����S-�y�K:��ؗ����G�p��J�Ɏ���d�$$�c
{3�[%����-��DA�L�o�Q=}���G���N�w��\0���d�hJ�5X<�=��t�.������,�dN�%�s'�5F��2���mtFJ_�3�W�&��[�Q������8��͝�v$#�`�{�w�ʈ�m�`���a¼9F4'�qt�����1�`�'�oJ`�'�e;ZY$���_�.�ǰ5��N�c�k����Z8j�S,�����D�yT����E�l�3q䋽9G���Y	��i$Z���Y��w�#;��9b���?����z��OM���
V�{=��j�40����.��@���;�}`��+g0:x:O�cF��O�B�e�80>�؊�τ�|JT���|���p<�̬�j���䊾�PI$�5~MV4��Ὤ�~"���{����
�R��C��v�4�9�l_�q��/[��� 3:���K�_����R2�;M�K䃫��g�7��7}��:on��G��di�jcU0�|�Ű�{K�ֺ���A��*Fnc=��s�*��.Ԉ�G?���	��Z2��̭��<���6�.�v^�)4�9��sH�pׇ������J-�aĆ����_�Dg
�]'w�M��H9s�{f�m�F�3{~��5R�������s���r)-��~T�b.,�a��#$'R(�kԈ	��o�4v�	�җ!0Q��� X�Q>a"�Z�WNn���tIf���$*S�4�/`G�e�l���	�m�RMz%Ͼ�I��m�?�� �4��n�����^��8��βMA� ���7�e
j��)��r��Jj)�Q��m��鈑�����a��jg�c�kP��Eׄ$�<��!��[uj�?�T*~wN3�|s˴ c
a֔���<wB�XS����a>^L��pf2o����ܵ��.���K�����Q�s�;2��`�`�����1���AS��V�=��#^G�3娄W�}��jb5�[f�\�$:C��/#/�>�ñAH xFn�FH��$�@�𙚀��ݙ0��R�؛ D��<l�_�7E� 7-�U�nRX⠈�XŌAV�@gIZnj�=�p%1<̶�W�^
(�uIB��!����5���8�j6a��
�ʓ�Jd�G[��*�QP�>�X�n����To�`!���n	�u��5оj���*m���2��/���b\�S3�� �y��J�'�d�7݄�C��y�&p���G��FTy=�~��X��R��s��;q三{Ԃ���}Oҫ����0 ���L,����o^��tS�4��:��#��~��M�¦Fޑ�6�<dT�pi�S�#X��6��ϧ�vp�gI��B_���_�E���9�I���)#�[��L�,r7���ar�D|��mv���"�2�!f�G��[��#g��+	�����7����w�d�~2�Tj�s���a=j�,fڢ������S	l�%�����XA |�1f�B.s�10]~Y�����5���vD���XA谙��h�~���Ǫ[?���;�K�E�P�iAE��9�ZcH�z��X���e�Ty���N f�B�z�y���8���\�dnq����M��j�� �נ;wn�	^���t���k�a��y'�O��������1,76���]3����Dh�PeW��m��/�Nd����q� ���ROUe���P2dx@�6"	xh�6�L'�Q²g�~�C\ I�2a��B��	QGt�Ꙫ'�a�G�5"Hs��e9i^mzޠ�p|�N`��p#��O��Xl�j��OⲼ�V����
]�m�E�/j�=��}"1�^�B��y.��v�\!�f��e�B*�R��Xq��s��Z!�~�E�;��Ё��TB ��x"៓3����e|D9�D�|\�M�Xߛ{]2�q��M�'.!�AE�/������'tUA�-,�c�t.B}���y╿��hǠC`���$�D��/���%�0#��Js��'�26�� ��=
.E�jt͔~s K[ r\ўL��)��Wν�TV���$d1����zԪ�bBٶ�ޓTg4=z��&^#L�HpD��@p(�}v��$����,����̚C�j���q��ޖ�� �Bk�[n�kФm��r��K��kr��ѷ���4\a����v���R��W��U;�"�w�N9�q�S�h�c���-ͳ{�JN�  ,J���Qp��0*�H��$�q<c��?�l����Mo��{�Lf�CI����� ���R��nxs|��D��˵���w}a��+��l7�a���܃*`��9�����,A�2��s������/�Н3 7<��^N�j�i��m��ڳD���~��$cK.Ʊc|�צ�>!���%�p����V-�ԣk��Yyh�hZ��.N��L�5�F�EW�=/�2f��y�Z-�4����!/��*�֟78���ʑ]dP4��k<V"3⁉��\��~$��**���;�{��a�6J�ԃ�07n��bkE���F/�6�-=��2��MU���=&���c��iϤs�BO�SvG�H�J\}Y7��uAn]�G1����ɄϦ��ᕅ�F�)^��5���������̞�̥>�X'����4� ����Q�_ez�C��]{�Z��{Y��ֶ5���u�e��{����
d����΍O���pW��00� ��fG��׍ ^��ߟ�-[�n�:P�G�	Y⊷ "��P�i����\�{�#:aB�F|�g�����4+��C��ţ��::f �&���C)��AN!�$oݐ�멨�N =��s'+L�}\ 3��z�*���A=,c�te�dV�� ��3��G�"��0ſ��q5��[�����TB*t�'�n2���x^�ś1z/a��/��������o�i���Tl<r ����ե-�w����I0^�W	��\#�LP����O�	��t�a(׬LlxNp�^Xe��v�gM�t���� F� n\A���Ud�d��۫��X�})��<��w�l���t=��Ġ�����_��Aؓ _7����S�{��,�~kh(x�N�MTs��m�,�3�5��X������(ò��c�� z;��)��_��aX�>n�xN0�M^B� ���?�Ү0�?WI~}�@A>���1���"�9�DZ/:@�B��1G2w5�pܣ1�K؊"`V���Y�9�EV���]�kF=|4p��d^��,�f�(�����fT1�+7=v�W��ļ�;a�W9���zr|�/4�W���,\Ҏ�@�x�ι�O����S?{U6����M���f���MgYX�I�W���ĺr&��Z�p}�ZL{��C"�Y�]BRS�(���Ccȶ���I˼���o$R�������1�}Ӌ@�d�ho5�ʜ���ڠ���� 5���j���@wG$#н�n������1J;�(C�	�S4o]/qme��nV�']6��*�3��mی�c�U %���&��b�_MZWX/�;�n�J�wk�/�~����%]�O6��I��{�v��5��'��1^�$2��kU�=@���I{랤@�M쥱ԯ߭_D���71�&�N"㒬�:���@I���*i}� ҮSJ3*��WɋH��Os�$ӈ+�"�YXű���YkۜǷ� T�I�������uj����o���ivD�4�'���̡�(1��S_7���;)$,������2�S%�1V�^��jɶ2c�v������7�����j���Oj(UO�*;�y�S�����!���������Ղ$W�]:�,B�,�W��u��L=��!��'�"Γ���_���U`�e;F%����\����j�o�g3s�}��Sd�<�6��nY?3#��Q�'d���8�V:�U�L�F���8a� �j�D�e$Bb�3��������ppi��ՓE�]�aV�kF�����HIcֆ����Q
֔^�k�]�@�s&�>�}k�si�t{:X��^��.�=����/�ܠ!�rsI�����h�\��\��&���~�Z�������"�%�����B\�����7(�%n����]��L*�#����.ڵR
v�y��g颣h�� �`$�Z!	�6+U�K֎�w��>f+���i�(����D'����{�D�-�����޲]}0Bj+;nZ��'V#[<��:SD]�a�l���(}B��Q�?	��ؠ��yKf|YC�?D�R��P���n^'�b��ْ��?�
��WY˄#Uy��B=���X,;ڠ~�]ww�~��ߵN���,0zrUˇdy�IM��'yƠ�9nȆic�%���^�`��}��r�➚���s3�U"�Q��J����ڮe4���%�}�簣6��lf��l�~0���3���;
��9 .�R�Fq2�C�w�n��_ ��x'�R$"u�#&hA��y-8�����u������#��4�+����*ɳ���G\��wz�Y�/�P��r�w軈��q�u��`N�ROx'�q?�Z	��k9d|;���:�Y%��LV�����7�:�^�ef�ʰ
�ʝ�8=ؒ�2��/����fx±n��d�R�IS0���@"��XP�A��8*r�d�{7k!�٩����Kǫ�=�[n��3a���V'�➞�zk�����D_9��̒M;��t:<����������7w�-A�#� QM��f��cv�^5����ϝ���,B�����ux�����QĚ�U���^��E��C����z*&��<��A]��9��/O-��p��[z_X��wX���In}�>ﳶ\;�L@�]H`R]��c��/���+�uI�-x��l��J�� �1�i�>�2�6F�՞F�\'���:�4�;�� �|����
!0�Y0p��ɮ�%)�Ɛn2���WR���s�A�c�����kD�1程f�e�	/�9�!�a�L
�W6�j�bHrB�`���0�*�I��9����Zc�������^�W���Ų��!K��$���p�Bzъ�uq�0�ӂ�BԢ�ʉ��BEq��"���J0~'��0�Q�E%δ�'�F'D;�{���KH��X��!���NV3�<�p˹q�v �c
�ht�y����������6T_��F��6���N�9rAF��Aa�*����J
ɣ?Ȉ�6O��su��"`q'oJ�.5&��l%i�Ճx�� b���;�yP#���#6��T7�.`n��3�hګ������rBw�U�������y �?N/K=�����m۩D�R�_������x���c�fX�s�I�ΥK��=kQ������5�%Os��9��u�ٮ��;��u�!��od�MӘ(��o��gVe�Ր\��a��ꊠ�r��ht�$��27h"���L0���:�E�0]KYn�@C_[����\F��E��q���L��dn�geݽq>$�G�;�	E�2�aS��}*K�%�V� ���c_��[���J��V-v�?�3W�:!cD���_��	�%��M�b3�J��ҦKZ�<���#�y�±v3��$�͙ϓ�'��5�o0��R;L7P��?��[G\�<W�M�.�g8�q��}�Moq'vW��T7��;22��k�B='n�e1l�{3)W�5�t�`���z��|�曗X�v%^��xμ�R��B���ɚ���N����s��ʋ�����;�2�ߖ��	]DEM<��+���b��E�;�Y{�����'d}r?1̔S>'m�U�Vڵ�M�'̦�?T�,���N���.�y�w�%)�ң�8�9,y�՘W
o'��`���^D6ws�� ģ~w�Xl�@����eA� c�)pE��z���x���oYr���vٽc��t\�7�>�`���b[P�-�TB�s��.��`ǭ.��,�rQ8
��$�y_�9�Sxn��H��v//�Nʶq7��F��^��S�{B=��Gᖔn���k 2?�� :�݇��v�7b�7����f��$�ֺƵ(!�c��qgC'#]:�e�"�;|���ı��K������`N�e�����}��܈F�_�T����)R����S����{�?N����7-6-:���� �v��P_���svx_�ٽ��z����G����lQ;`Z�=�$S�f5%��B�[-��g����2%�w�x��d5bO 1Oa�ߤ��'D�Ѥ�c��N`��4�5�B�l_�v���;�y��͓X5D/�z(�K.� ؒ���j�4��
+�g{`9���'n��s�����b�{|ϵf����S��;1�1� ˁ����ށ��$o9�C8���P����3�h�߫�f��ch��
c?)� �ү(]�����D�E�����	�L���1=���M�O�_�K��Ü����H����2�x�?�1�	�c��aˎO��$��q��!���O��H���L�0���.��u�(U�n���AE[�ɓ�f�������Cn���	%�	�)�W$���I@؜��� ?�����fy�o7!����or�3)�U�Q����B�d����A�Ń��8�;֤���ÒIRf&����u���x1O?�L�s���%�Dv�;Nj�@���Z�c!͉l��xq��l�q2ڋA욇4Y
t�cJ��9p��	�ػ�Z��  �z%B K������7h��Ƌ:tG,�Ef���2��~�/��r�)mOxJ)Yl 0�3��GOHcn5Ԛ�8��l���_e�X�v!	��s�R�)���a�m0U�X)���!J�+�=���3�"X�d��Zd@�7X�5���϶��fh�e�'�A��j�bO�霌-wm"���3�w�;0�:���a�������1��P��ܬ�
ݷ�1iv�����<F����7��뙝ɧ�������D"d'e���YE�y6w�Y;���8M�C��]��LSDk�X'����e{�u=Uf�_�\�.i�8��6�+��L���X�`dA�s�:��]�
�ֵhU
�I	=6��1u�̏�.Liœ��.xX����J� ��a}���H`'���55�9����x�.@�]��.E�g�
�ʇ�h,�<��:�.��V�bcR���=�"xgU��T.�#}����+ő4dZܟ�gA��ρ��~ՌGz��
�^�D����X���"��&4��L�-�)~[}J�~���WE�+)ਓ�3k7��*�ew~�?b�ط��ݍ��$�����it�+l��@�YD��c�_ؠ���e Q+�'�����MY���OȤr��_�Y�p{t ���]߀x����^��}z�*��A��D�s,�����o$�Ź��~��Tg2WZ4a<yeu��ŵ0*V�G�t�Qs����N�}�b/������tʢV����e����KJf��/�F��4�wr���w�cA��o}:�^$�SY�X��9�3y���<{F�eF�6�������� ��)H�UJ3S���5�{>n<�Y�"�drX3�l�|P�Q���Fj�qI�2�p����b�2kg#�����יq0h� ;��
�p�z?�JX�'�H�0��X7����=3�٩e�f�&�'���`
8.��i1%���j��/2�Z �Xz�e&����+^Qd-�@y-N�	jb���;��ͭ#ө���ebb�f��Q�0� �i���4K^�.m>N����8�t?뚎*�D�3p;��H�L���O~Q09{�I]��8�[�?��)��.ddǨ[uF6D\3�oi�.A�K�)���7����u��[K�Q�d�sc*����z���8;�����/*c��e��z�xұ{n��e�M�P�����i�_2^�S38��uN�_��Wv�7��� ߋSS�>��Zy�i�-��+Z�g�����$i?�b'�/q�K����c�v���B�`��	���ԧ�S�B�Y}\~����娳VH٩"���[���������)��\�vxK�-��}�.K��ٽ�`#�%�@�4�8�Y*���`��e*���63m?mʂI��Ͻ�V"��,���sO$�!D��G/Y�.�K�I�<��a�$���z�rh�G>��g=}�>gd�ū�R4�g: �{��|�}a)ue�Z�����${
�2����� �	h�Ȗ�<�n�� N%�O^b��{��+��VǕ�?_�,l
�d���+T��c��&j�����6�3�M���˝?�b��mp&�6�vۓ>�~r�~}C(U���,0�b�ch#=r�����u�e �*4j��dT�.��|t��t9g�D�>G��M���t��P<��.u���/ETl����(18<�#w{\�*�R�N{K�7	��wn;A��ݨݻ�m�O��`��X�Hh�����H���:w� ��2���n������0��ꁃ�	 ����5�QX���^�cK�����'�$v�$�����&��W����K�&�^ 	r�ݻ�3���y�L*N)L�X������}�N.�!ʕ�A��`*`���lQ��/�e�+)ͭ�����l�=�?�x �m*��+y1�p�l�7l���`���,����/C%D�;6}"sdY��ixU�.��
S�bј���C�0��{��/	oe�F@���+��L����l�t�t���T%$G��q�F����ER0��t8t�"�Ȼs=T�|���x���o{<���%WS�҃�R���";���%�-���f�������g�՟.� �-�=�0?_;pn*Z�?���k�T��2�����I�x ?(UԢ����$Bq�?|� _�DsJr��F��j���^~��Ů�'9�D�^Ԏ��J���� ��9/L�ĪΜ�2��X�@[��S8q���ln�`K�R������v�C���W� J.����b�d�R�X�����{���#ϳ\���ٝ�!���1��y���]�ݲer�7&�QY23�Fc��D��a0^�9���)��.'I�[#yK����*�ǰ4�H?�V��i6~88eԚ{t�v���;F�d�}�BYq�.'���{/"�aZ�=b���Q�p���mnf�Hs�uJ������JɇPF3}�@C~��9Bh�J�:�S�6+�I�V��h�܉:�ߧ��t������ɰW)a���T��c�g�"`Pqҥ����9�h�v~)�\k��Fcba:����
P�|�1�{N����,�2��.��6�5FP���a�O#"t�F�@ ������5����Z��ʋ��??[��yGG�$���K�b���jҎ��dD���:j�a(*��8h��]�P�h*9��o���-O�&���h���G�z�$��Hmw���Y��L�\��k�� ��,����k�4.�sm2�C	5G�ݽb��1��gI�T?�*�����m� :tv�g��o�����9�߂����Ǭ�|��t���@sh����i
��Ve8)�ޯ@�!qŻ����"�&�2�����UvC���� �:���=P+XzG�H��3��xmp]މF�ރ/7��{<c�h��7h�P�X����B�?�3�н�O	o�	f���d<�����0�R�&���-x��9+m�@> ���lRW���$�����=@73݇��������ug,%됿j�Qݩk2�
hت(����CG$
X K&���¶����U�\	�C��<�S��f�Ⱦ�hp(�^�k��lX-ܙ�l���-+
��"�0�"�:,�G?eIy����
l�ND0��]mP�g���bq!�>�t$O�^fovjǷxKC��X
����;z�)h�λ�c�|�iXX��I3���8U�Rك���#A��OxґLìЭ�͘����Y=�U�H�&5biJ�/(h.�G2aQow;�����@��G�	
(�����s�s��_͢�mu�u/�S��͌N-'�U�s�k��Ç�C3�� 8�O�:aNL����?2��e2
��.���At��d
�4-���e�[3RU�ȏ��9��ߛ*��跇ô�-;�i�Kܮ ŵ�Jk_�h߇�;�������)�+��`��i��A�P�v�'t��>�Ƹ�.;Q1 ~���}iR���P+@WX7T��4-�J']�_�0H�%�-9�x�E��jH.l6Je�^�N��F�����|���]�ͣY��Il�3jX׭E�3T<�B׵�)��qzq��V��}�m$͟�xO-Q���M���e/e�#��ѨJ4>��t�]���	�v$��;�2�'���S�9e;��I81����O�[�>��F{�D;�����DT&��iRlqa�%�k�K�a��\�/�45�q
�buo��Tge����;Vi��XE�5�(��\�&.�Ӫ�1���~�����*z޹Ո���)���Ǳ�9�Xu,����\��b	=��_�U-�Y�'��r	����c*�ē0W�sbV- �N��-�2z<���Po��K#_xE����à?�|��Q�a_n}��LW�qz׾�����[��ٌS��z���z���j^����P�S>����x�u�#�`��\}j^�Da���x�E��>�8�r�y��[��yZ
bk:������Vtz�P	�8q�`��:���ѫ㌈Y��P�4:9;7r�Նy۱���A���R:^�����-:�Y�)�H�K@�3�&W:�Xf����=	>����M#=��S��N�?����Ĉ�|Pw���f��\zbw�z��t7�=&5���-hT�ʧݞ�D�O�oPA	�_�A�bv�[�9a�g/�Mj����>,f���W���	�a�$gL� �IoudNQ�Ӽxy��=�1�*�m<��e��+w�*-��kK� .���ePU&�w鶪O7nG<�s�
1��/A�Z�m[ܗd�{�Jֺ����?�H?��5j��G��.o��p����&�?F��o j{m�ͨbC��9ʽg:�
�N[*�?���vH�wz��t���bT�EU5[x��~��Wߩ��<�l��!����y'U'K��LAz�6*Z���2@)�y�;���B��HԆ�!���쬿���(o����Ƶn2`�a��� kf?�� ү��9jQ�l:�H	���db��b0�B%��R��xF~����J�w���(e��(
��Oc�»H̎�g�:���\f������7x�����]E^M��ى�yn��3�A�TIp۴�w�^�rS�[��{��ׯ8YW?��jZ&��н��G����E�!_%rϿ*5*W_������]_��u2oN��2fKU�_��@�Շ���ön��e�l�@�� /!#/�LD��O���^�A���V$��NŚ�$N��r��$	lӱ�H���Y�(TJ�^���I9í�?�^5�p�Կ=���:�(]��^V��]}-RV���G�q�)��}��nm\�a��{X9�c�g����Q�w@<�lϩ�Y�uT�`5	y]h���`Y&9���.����GD�l^=�mqs�zX ���w��N�
�f5#�3�k�*J�E�3��>�6�����`/�x+>�p򦦇��|�T�T�G�sg�~�#.Yvf�$0a��Jíz��Z":�'���%�8>���T�:�Y�H��˓��D:�e�/{��"oU;Q��2+^EKTURa��VT�h��W�ϓ�(AsM��+Elԩ�	b�ZɌ�`���ħl�Qw���<+zk��)�=k;ز�{o�k�h��v%�e�{(��)������iۏ5<�rŃt��]�a�o�Y!q�����ʂb9��̴2�l����j!:�%s�����f��X��9���} �.O'3�oN8o2�aK�PE�o�HE�l�GA�/�I�)L�ت�	�ΰ�I�Ь�_��~C��NP:�{8�#���,��n>؟u�n�#*�~���u@pq�L������ܘЮ\�&����@�2K/v�}��&iwE+H�nm�SJ�pL��/�avH�,��k�*^ȅ����	0<�6d�NP�F������b��~�?R�� j���L�ϕ���ya[�8^��V`�&ւ�=�ZS��ӭج6OrNw���!׬P�Xk&��g��hH�7er��a��_)<�.dO:����-��o�%,�`ŏ��k�b��e��E��R*Vcc-�����@�D��#��uk�k~ YO�����z\����U�y�����|���%j�r]��(��=hE1�M�9�\%zh��������d4ѾT!���?nNN-�%1%/`�i��Bw���K��-����lx�^~��yǓ��a�ғ��{%���i�?�V�g���N�i�	�k�0 �='yޮ8��C��9��;��s��Nt�[�Ƙĩ����'Hw�~�Ċ}�K�n%��\<��U���9ϡ�ͼ���؜����?5j��^,w8���~�?'zr4+댯�+]���[��_~G��(��g�ܦ� �Q��]ǝ��4��(��~&�H�V%�� ��.�XP����71���ӌ���(�a��?&�2�kK��wU�X]<jY��*bx'#yU_�5���|�PS4�Ն������8�qm ��}ƝB�/�_�M��i�d��P��ߗ�8�Bk�yچ\�Sh?��AG�|d Mf/�+2�t�'�I|9�:�M���&wl6G�<��y@npC
�k��t�ު�,� ��%��'��e!L7�%̊����"M�<tN�X�=�u��ńx�ι��ĉՀ~�4n��2?!v�=�B2�JE0EJ�`z~�c2�U�R�(�*�����=-V�u$��7���Am��Dar�(,໶j��tg+)]�f?���8.	���:TF�-�wȟ�������UO��`��2��>��
�?`,��|  �L��]]s{�[��sz�ϽW�}(D�0S���I��>�k�I��2%�/���8K���b()����z�ˮ"�j\,gI���a���ݥ��龊*�}�����5�M%����j�ǧ�uz+n,�9��f�>�m��U��ʱ��R(m��U2�Z�����6$4����C٥��̬��G�솭`z^ԆnI�Ϧ�6; �Y_FS�_�3����'���m��w�.��ԋⱣ���S?b�@���݆����;�_7�L��"x�[p�1� �"���p���������Ɨ���{�Q	�.�7���ݢ�W��.��\��O�Я�QKoZ�E[}��e
���>��v]�g��_���f�ч��sy�0V��ݍ�A���ͣ\�y����(g���6(�i���D~۝����1��,�F����,�)&1�XҼ'8�ƅZ9A�<�q�L1P�����.h���[�1\��J�-�/�����J�"�/bGnd>�5 ���c�����C���"j*m'���*�N�>]��,�?�*l?nZvz)d���rht*FWCð �<����)ΓO߶��w.�.����'�a}NL~�|�i[��_F�,���z&KI&],G�B����ΤE��:e}a pd��A��:H��
���4��
��I/㔃)gc�/�(O�G�E�֝���{�He�ֿ
a� o�o���tr���J�Q���o�E6)�\B<i�	��G�@eq�͙M�\�z�Խd��{�DQ��as�q]�´V�F���x/Z�d쭘:@G�2�^���ڂ�Uo���towS���͠��/$��A֛�_��O���ǀ�=�ZR@��0x���js�m�����g=֏��q�g�CWj���uAK	[Ze�7�*txKw��L�c�L1�vw�����g:�3Z	��������)6}�2Ц��Z��RN�r=���:ʉR�t|Sӎ�����3��;"w�P]�?���1���_>DW�����ɄW�;C�8���y�/G��]�X.�(y^�G'����Q\���2Ò��޻����<�pү�|d�
Fj���	Y��Vr)�L� ��9��g��� �,$���)$e���FdzX}����,%\]}��s�N�4-,Ց���&-�[�0���.My�
K��2V���"(N6�b��e��H6���� �g+���Yy��E�ȸ�y`�ѫ?�S�XNSAh�	:>Z�v�(�"US�'��CM��>�m�����уE =^A����4�B�Ȋ�f����)�1�6b����M�l�[
�}�H'V��x�=�vw�D�c���(��f	Q�����]&�Cf���Z��T�bb�3�腫�jlt/�Mf;�c	��>�㹯�*q�JHQ�j�W ��ke?��{aV/b � ��p��Y��]�.��P#�������*��-���&,��,p��k�V�pQ�A�m�qڇh7-��N������9����c�*a��B��1�t�!�:䷎��bz���dU�MXb*�2X�������\�+D+˕l\� ��9�N���K���
��o���Ƌ��{���<�t/,����m$�@��Vۻna.��	>I(2+)1�e�јv����ƺ�7+���S7ٻo�N�NDw)8���u�~�.V�V&�E�'���^'���E��\����@hd<!T��f��|��b	���A.2Y5�}���(@<%;��fP�?WF�Ll�������S����-�s�>�]t����scą��f���C����#��������@��-Dj��R�J}���a����"����(AxH�*�1(�X� �ߍH�ٝԃ����ݘ��mg�i���Yx��l3����X�����:�4@�O1�L%y�ֈ�H[ۓp�L8�T�s豌i�)%q�����{Dq�3d���(,J��G�h-s�P��;I�z�鹇>�gM֗~�^�w�^G{��*<=s�&V I(�M��ǣ���"�vWB!��j뎙�q�G%v&��#��T����q&b��>���4���x����*��m)�O���!B�9����t�t8�<����ޙȑ/��|���E�Y2����ӝ�:i�Pk�6O(^H��4A�����~p�l��c���"�\��e�*�[�(]��
��;~�� �O�s:�h?	D�C�G�H�ó����յ�ƕ��*���x�y��%�%|���9p��Et��� �:��|6�(~�&�R�Qo7�����9�A���{�V/`��<�e�h6����ң����t��6��u�Dv�Uڀ�7jɞ�'���>*j�2���8(�6j���x{)�H�<h��o2�y���K�Y���9��(��-ģU�(l���w @xb�Ϥ�a��ΎJ8���d��t�#���D���ߴ�'щ�r)�[�b������(3G惻a`\9����t�����Y.��()u���B	���(@]���	�߬�H��řs�/X-�yU�����Ա���P�=L����M��ƙ��~�k`ʝ��Y��������{B��Ij�h�$b��^�WT�H��@���X��ͧC��e�Ԯq�#.";�驱R�*���i� ���~�f5+��� &�U��>�4v��ȉl�Q�Ù��E���ד�|�ɹ-�����AGxj�Q��K�����Ts:�0�x�L(�v�b���H[�M:V����-jY;��Fm����u�Ș}bL>���~w8(�/�H�-M$�ԱZs%P�7�:ގ�?E������s��vxU2�`Ē�锅���l�$�ɂ�H	�6'r�	�R�EA!b�f��
�ve�C���e�Xw5��ﰽ�%I���a�A��W:К,!�9IH������&A<zjZ���it���s���f�U���,O=@��)92Cv�4��\hC-(�cu��Ldk]���ml�b#�`�D��ف/����S���}|���gJR�EP��򺵮j�#�֘�W�`x�?��
m:NG�A74Ja�G�+���w��]�����~�@i9��w���k?���0�VH���>��*MÕ5�7	�'��c?-�ec�tt��2|��u8�tU)��'����3��R��9A�R\S�A���b��"2@���n�Z�����{UR_\�y�"k�k�屈����9:1�=�fb�>����A��:R�S�#*�@4P�L7����z�vsj����d���丫�?�{qB�f+��9���l�IU&�J[�{�F��D?��nNz�uk2x�\H�h�@�0�	��eխR��)eI=Oi!c#@�c� ���� ̄ޛ�S��������^N��`3�R��'�c=�'�J����J<ȴu���!a*
�r`��Er$3�������^���NIi?�BO�#�sA�N���vt&]��Л�E��v��R$$��!ϐ��=���D� K�I���r������[�f��IG	��������d*R��f�x��P���r�̝Z׶���H~�����]Ѓʊͨ���˄�����ਉ���a���I��7,`7�F�N����"�L�K1l]��7�Cy�`�QH�d2�Ip��{hhhV(�4̟��,�Xi�y�e�l�g� ��%�`>e(%��~u����gԡ`��6)%���YĢ`�נ�Ωʫ,�מ���}*������0=���N��8.�q�����}8��U����e۱@���V8��y�K��w�b��|�?V,R��x���)� ebw�C���݄E~�Xͬ�ùȐZF�iFZg��^Ð:E]1b�K{*vP��Z�Xs��]�dG��p�=5��ǁ&�d� �	w�{,r���#�61өO�+LH�Ig#�- ��h��|:��WA�7z����*qϒ�D���'�v������"�{�����f{��c���4�[F�Tj�Y�͋ި
�T�g�L 5`�0X־�I��∂�)��l�;.�D�=��A/�'�\�.%��`x:�[�W�m$���3n��O~�p����\�׍��M��tTD`�v�O����I�Q~�և8��bP�ڸe�h�/��{�	u�eK��ci!@���`�1���T[����o�\>A�㔖�A�Wi o�j�N=@5H�K0ְ�8�S�=���_�cU���^{���Vojm�¼;����.��s���w?�\jB��6��|�a3�y�yF���5CŚ���H�"PX2����D<��~���	�B�q�JÚ?r��T"��g�*�m*	��%�1��qY��P�TJL������'ש=�9/zI_�v���X���\��:�z���fr����8��������+��\H��f�>hh�(k#�N�t`v��$�ERb ��@����J ���f�HJ�͵�& F����:��m!�¬�P����EM���}�pW�I��%g]�9���fT0 �}��Žw��h��<QQ�Ǫ>���P����G\B �f�uӧ#�;���6�ePq����Ϸ>�i�z?�'f�����Y�~̨�э�.拰���Z���k�a����	�?���d���)B�4�E�;��b[��Мve�u�Q��<��/3Q8xƄ�M%[�7aq򵕷,�ݸޓ�|�'_�ݻ��7�ŋc���4��7y��u�O e��V�=q',��Z������'���9ڵ7 �!!���;�x�V�X�BZ��0xH�B�+T�C����2!�n*�4����*��:6�v�����l1����G�З8};��t� ���C*r�֭�!r�� B�}S�Ri����~$tj}@�}=�e5l�X�yN���5��l���r���sėli��-��5 �a�z[*��F�1� �ŝ��ImaMW��ew��9Pû7�~l�e�-�J�k�&�/z�B=�� ����)]9�M�@���cx[��1�%�]f�?7te��[<��ɩ0>�~+�8b$�(�ǲuK&g��EJѭHgf�?� �m�����Ú�ӎ�{#�E.�P�Sy� �Xp�]���Ҏ��ЖtH��JO�ܤ~�(ƀ�$Qbg���6װ�sIXx+Z�G~��B�Y�!oз}`�?�f�KxӠ��g �}�M@�H�sB���Q�T4d���)��u`~��О�����У
���0�����l�}�<���A���HT��m��,� ��ȻE�)�c��]V��d;��߽�F`I\'�-}X��o=�Κ�!)u#U�;/��ִލ=��M�Ϻ��h�DL�e����������z}kc��LWz3EuMU/��8�uW��v��w�%F���j;�-68���f�qPop>L��V��C�1%�r�������F����R1� ��4Nf��@_�5D�q��-%n@�S�r����C����g���ȟd�Cho{��y��=S}�F�u��l�P4ƚ!�x�C :�I;�Y�h�|���{N���pJ�i�����Q
���-9ƽP���o�}��GT���CM(�\�zq��ex��������A�oS�~6Pp�~}��t'�����f�^GB�)0���/���Ǫ�<E9�Ҷ������
>۟�0?I�!h-!�����\NbH�v�M�hF�`j�2iju�]-g�9�Z��l��?��i�!��lxW͢:#��k�C�
�%}e��!�FUo#�Zt�)$�g�������&�u���+W�Al���	z|`:��}$�+��I+H	ͱ޽5��1X��)|�j���
c2�O[�٘JGIv��Zձ1`��Zb�*�����d�Kau(<����xH���J���g��(�Wtݔu�#�k����a`�\��C���B7�p4hM�Yq��;�s��#2��E�[�6�p�=��a�փVy�磍Z��^��i���@B&�L��RMuWՏݿg] \�Mß��\������>���< @�?k��7��x�b��)�x}������ֶ�������*�.��v;Oz�@�{z����P�جB�i$'m����WL��Z�o&����~��-������?:����7R����m>�oQV�G�ꘉ���o�m��,����bJ���&�/Km(w��H�.�c�P/�Ά���e�|E�h��)q�|��/��]|e����0��&�.�x�N���!��0Q*����5�}1z��*H���l������|��@��gi�Wh��D����Qm�U=r���~�9/	_�O�1NoS��i]�g�~�!�6��mQ��】��o�h��dSp�K�fy,���<!�RZ�-?��<��cF���X�7_1��?�R'j�Mú2Q������l��&�9`j�~st�rɄ�|�T�=����B=q��8*�����M���9� J�Z��N0�C�þKN��aC&�To�(�u�B����M��$�M$oQ�C��K�tt��(�Bg�>��`%B��D��s��4�_�Y�<�|i����e)`�*<�&���̟�h�����/aP��&d���.�H��fj�<lC�-�g�Մ55������J9w� ��[u����Y��$��x���6�y�l�� ~�Ǯ��٫��)0��]��Fq��O+'�O�-�|ߥ)���}�a��_�_Q��C=��-Ɗ6�)�����/�8nx5��A��i��ʌ��(�7��kf�Ԛ�����,p�R;�'���;F��"���r�gp���k�7
;A��t.`c�ň�p���
EU�ͧ������뉥k�����ʬơ���;�M�dCW�]@�f�&k�"���<���f�X7<]4�yz�����G^(5�A�-E�p�,�;���qyDP�BM�f�8�/|����q*-�\�˃(G ߖ%Ǩ�����u H̄�-*�}d����y]�l:"Q�͏vaY3܋}۴����*\��q�
"��&/��?���i��y�ZX�ޑ��L�I}Z?ZI� :���ʓ�c�s�Ҵ�mh�����K�QA�����4E �w r���tN�T����U���D����{#\�"��t�m-�I�����t�m�w�eL���w+Ub8H�w��6W��&�ܶM&��~��G�ׂ��R����z�D-١�cH����6(�y[1���H��5��M%}�T�c���2���V�8�g����n��@r!�f��.��'�a5�\���\��p��?��'љG���B�b��Wb@3i�d'0���zЈ-�吊�f�N����U��-��Zw^|��ī�>�%-���X���p��/��^�)�74��4�!"�uF�`�9��,����f����j|����ZV7Mf�$�e/�+R��>�6��6�����'D��ʹR�J��o���Ox�qgh�����-���΋77�$k����%�����B�N��#=���$��9�j-U�Q�<�-W�q^-��&w*���}��3^�Z+}�!L"2��5�:%�S�޲�����WثRt����Bi:eԊX��Q���� hx[�[i�)�~Q��6H����9��N<X�Y�#�uk�S�y�lq7Q��{PtܳI�,&�S�*��E��$F�nNE�x4�lWyu�ݹ�a���W���K+<f�m�}�2�{Y��Ys	��r�{&	���|Wl��l�U93+p�H~ԣO��w`d=o�Z��*�6��C瞣v֥���0*x�1*��%�E��,��1�"�U ��%��"5�e���$�L� �V�O0J�HLA�����S�ػ𢯄��o~�̒�2"@�h�~]��?�Q�w��nu-�1�B�ی� y%`c������:�S�h/��g���}C��<(�_.9z���p����U����蓞E��a�S���q��3��<�v�Li�n	g�%���|ty�ɪ�XF�8�5����h~r"])M�+���I1���>� :��K��d��6��p4�N�0��8%�]Nx�fN��יg�V���R=�k'd*�e�l�Pc_Oq ރ�#(G�wM�.l�����ӥ �UCkw���%�\�T�J���p� -��@t�y�����=�¡��`��!2�kxB1��t7�D���TaDλ�y�g�>O19�d��	�y,9��K&�S?�2��OK�pʶ���#Ö#�sr3�Os�������$_�M] 0����aX`KjBWh�� {�0e��u4.3�0ݖ[ִ����� 	��v�VǒL�ɹ������|���P�Y��q�p9��@��@�n@���0��b�3�C��rY�`M)����@��4rr�[�.��j������n#h���ށ0pǁCT7�ʙ�=��G^�<�ŏ
Mx�671�3oOe���䵬9�D|/,�m����ȹ��M뙨��'�Iz�5|�>W��:BI0�������>ْUq���dH_9�����4E����o^�](ֲ(G�Ƣ.,��7��d֑\o�g���pd<��r7	N1�\�H�Ye�)+�p,��q֔�&�O��(�в����jM�T`A�;FHh�N���-4j*H���=����/���0J@a������"&H���)ť�׉F���q;W���iF�ԻSOfO��B~7,1��/���5s���~`8����w���c�Ge�f��ltG�dZ��3�|5�6���I�pJ�3��_�+|w/��i|lާ�	�G������ಆo�٠�S������h�H�BUDW��u�ul�^�C��,��]�\F|�0��A��:zoY�1
L��Y���Y�DK��]��V�p�_���� �BIB������2ߝ(��N���^Ow��Ӯ�i"�J�+郐/����i���ڬ��d�馁Z���I� ��{�!$�db�j�Q�ǐ�?���Z�3���Ezȹ�>˄n�aF찃2���"a��""D�ǔ+�X��k̈�5 �"~ܜ�^���~'X��C�
�F����?A�[E�A7�!A��0Au����v,Af2��e����rT�����`%<�����^M�����������vL�z��#3K�w�]�B<~ �
��uw������8f���e��*�����A��V�@�^�c���8}��#��H�E���:E�z:<����� ���#C��U�S�4E��[+¦_Oi~��bl�Q%��_�����>��;���R{�L��8�rb�wѱ@�"Lj�OTK��L�{���ie�(�u�s|�R���ֿE%bb���mq���Qv���O<u/S����f�a��8}�w�	��<Yƪ��L����'ӽ*��Ӧ�\0iW�mg�M@��\��҄!ƞ{l��E�͠���};���?�]t@�ɼ�%�h�sX��w�iuIeB���ThX=k��� ����/��?m�z��a6��~��V�ѻH�F�y�@{Ve���ZƖ���ޖ���C����4�� 3Օ�'Z����C���c�C1��W:���T��¥��[����;�.H��tw�=��uJ��	@m:!��¤oᇊ/@U�g��\��Sſ�*`I�&Em~8�*��=V�^������.�hrˋ�I�4kcƅ)��q"+�ڀ�+���9p�Yƙ���&�
�ƇF�7�ܝ����#ٿ�7�*��ɍ�\6��S2������J�]81W�S�9�.i��W��%$X�Y���4�H�B��[ �C�UK6�Ԡ�dV����ͽ�~��
T;�ey�]�^ػ؄RhDEv�X��}���x�P�*R�*N��o �ನ��L9L�X|Ό����=���e�|����
��(�>1���rH$]pU���G��G���9-W�宐5�����c���>b\Ri?P��1Y�<�V�E�q����t�Kv�<��ջ���@��т�~S�
Ca/���7c���Nu�e(�L������N���}��L��NG�����S����rޮ���MRc\U��l>����P�H�*r�b���S�S>]09YˡS#^J����Ut���Q �yuW���������9E?��X)��'��[{�'���l>��d�ҵq��T�/�a��VO�w�;4~ij�.B��82�R������1 	4�>�q��8y�<坉+��Ӹf���˽�Qd{�s&=���=D�+Ѳu��v�{�H�� &Z�y�����!dcT�_h1ԟᵇA%^�"C����^xo:J6/�E�QX1}��7ѐ.���*�����U ����^�'ͫ����+��C#ofsL3�?_�5�QB��g�$
{v}s�����6���� 3���^3%L%����N��I�'p��@6�A�d��@l��J� r$����0�Y��%}�N��0q	}I����	o�x�{֖�2�1�tN&C��!7��Q* ��)�D�a���"x��Ƭsք�X|��\�U���?.Q�|�H�wB��e�.�� �Ulp��qphf�,�^�ǹJP3,^�Ғfa�Jf�p���z��¥�x9`��
��/�p�ډ6��QFщfi�L�XYfe���^�QU>"�����q&�i�����jAV�̹5��%����K���O�����z�Q���]���F�lQp����k�ìT+���#�{�5�/���
�l����sLѡ�	(^ie�Q�������Q�;O�W׀�Wː�h�G�C��#�B�M�4����L�+̊�r���Lu�a�:�+����z9�w.f��������	�,�&�=C��[�f@|��pA���`U	bF���N(��/�[���!8��L��(6��Ŏ?��P��g�{��M_c�5���c�/%t��w3�=�qZl,�1��4Pă��QS��i��'R�����y���� 2�knt)�OV\�D�u�-�L�w��r��_��BD~�45ɢ����m��b��t|x�+ ^ �7�sn�~��䤑�"n���h���F���4����~4q��~�*6�_������闅t3�08��� F5S5D�n�B�O��$OmȔ�M�C���Ú�d�Q�2Y*R��+���� w��&!b��Vu:���p�~��LT�z��x���/Y��� ��)���=��A��.2��� �Q�wt�[n	�T��e��Xd�L�Eµx}��!u��en|k���2�	ɠ-�-��1���S������0|����f�!��&�y����?/7o8q8d�YC�K3����Vr�Y��8p	$9��8�D|��q?�\b�Ѡ\�hjI�͇_Ym�:���5V(�'�Đ��4O7�?l44IL�Ξz�u�1���5� ���Z>�,R ��ǤV�c=�f�8�?pO����96Qm��`-Н%i���d�Eʯ[{�9U`��o�xG���i5��U�ړ��1^�LH��Wp�.7g��VL��؍��u�U���=3Z?�|yݷ�0�s� L|7q�A rw�Om5�>o�=�z[E�M����O��o�^�����В�`͏�P��t�^zjs�.���'g�&�̓Q<Vܚ�*Nz<7��\�]zU;uq�쁏U�̢0K��-��z�d��Z��b�v���[�vpS�r%="�'�0g\/��^A�y�u������#MX1�������2T��8���lT��R-7ʜ�����[�:`/���g�:����r�W!3�V�T1P�q+�WF<µ���P�t%c���&�>�����p�I�5 7���2:\��֌nvbu��IR53��Z�w�7n�0����!��n��~]$� ��=#G��lc#�F@I֪���cǠX�(u`E���X��$wn5��b�͸�r�{�oL��[�Ő���wM���)*����gnr�͞6���s��u����ۇ�����d�����f|�����Q΀���{���پ�=�Z��f~AO���?��ψ�������)�dZK���#术f��9**p�|���?��m}���#��l����eK^��ꏃ�V��: �=
�MZ�җ*/�EB�wW��G'Uר����zy�ј���� z�կp�+�py��޼!�dZz�J����7ւ?v�������!Տn��in
Av�`r[�F���$��a���w��iq`��$y�q��T[y��� d8sv4-�A}C+�Óc�kO��%:|_'ށئ`B����������BK��Vh����D��`��㪘�x�7R��3��RJ���`<��.�dPT ��\p�[KT��%��8����V�x��aP�ď�:"������6��w�6I1B���Ahp���0��Vs�Dir�
C)�a@�C�c/l�����z�me�L�J��|}��[��#-�j��������"���##����x�j�=��_�7(��2�q۰��`�C�1�n��U�$k�t������٬����ض�%�i�c�����ym筴mu��W3P׎d�\���6�J�B�����њ۝r"F�.�r`��D>D�G����^,x�|���]B��:�T]s1�B�����ʬ1���dUM�簼0� _܏[�b�\�dg����֮W�z/��q�9��\��˞�!�ӏI��+�'�ǪlG��J<j%B��\+����Y�4����B�v�K�1ʣw���ڤ"0�#[�F ���\!�3.La�4t3:��t_�TmM�<*�T��fT�V�I�S9eZu`=Qv�h�=GP�#�M�!��Ƶ2�	�����2�sf,��-:S@�z�Y��(\U_�b�h��݉4��>c��Y@�5�mU�W'��غ4��p�(H����eP��+�ي�*S�7Ձ�ewX��K�@+j5��P�{
ʈTfȞÆ��S���5�����'���a�5�QE=|�鿲�݇X�2CT��e�����z���O�h�GNTӲD
a��#�g�S�@�O�ӯ���DV�- �0�@��e�/�J���J�"�l��ekS���C}����W5���v�Q�K� ��^[���w����glO�ͱ�mW�>�0H��N(@�5��|u��(�u�C/�����h·��HΧ|Y/;�5���Կ�	P��p3��Ǳ�]�o{�Hz<�u}W϶<M�0L�K����8BK( 
%γW���P���өXS�����9첝��@%7���D�xMs���é�ʹ�pQ���f�$�ο�ًf�I�UiNȐp�Ϥ2���YdE����D�i�sd�v��ȇ��'�V[�Y#<����!}o%v@	�E{\K��0�i,��dY�*U��+BϊfmjUQ�m_���}��c/�7XIb﹟D�XX�#��$�߲H\Z��p��8��Z�=Y#���#��U~Ř���"�TNB}�\b���-b�'&���4��6�U��0R�[�E����J�/	 J1���_���r��������`<e�ݮ�ĉȳ"���#��0�D�p	J�,���C �G���yf����6.��QX ;��̴�9T�E�(��YyQ��S��v:0���~j'�~e�vZ�ϐ�gl�j7(�T�$�<�L.�$rڟñ��%`���*���z����b��9�d���{"��^`����3٣��'��ЈhVwo/(Ǖ�5[�]���c�E҆�<j]��P�������m))O�ע����P�&m�X�(R�BM)��H}�M��Ub�M��5�e;��NL��)�q�&��[�1ݧcjQ����Ke�!�=)�l��-�7�:9����Ám��I������F�~��H`~�AGr�M)J�ӯ>��te�Vx1ǜ�Co��8���ϔ��$�1mh�̧p�t/&]����H�h��`�H![ߟ�	��@�!ς�ށ�.��$��%�XSȑ`='�&	�jCf�\4��:K)�}�kC��Ƕ�$L֓A��s������t <{FZ�Իt���?�N/(6E�9߫�Bw��� *����Z�s�E�B����ֹi����A$#�c�?��jm�چع�<u�j���ؑ�㐎	a�	�=�᝼�S��F����@3���y����_��l}���C;s�7S�1���ì��6��$�s
WO�I�PG����'T��E�a[�.d���b�\jC|��F���{���V���t�'(m�n�	1@��,{�a~8�0b������t,h�X��I09h�Fvp�d�5�(���ъ�tz���5I�(v-��L&a}�3�#�Tgd����F<-���=,X��[��L���r4x��Z���.�����p��������N�V �@�o3���ҏH@�M�?��]dF�p�1��F�����t�d�NN�I֌���ak�1 �E@�"��z�<ޡӎo�-YA	�~b��nm'uH�����\��~��.�h��R�B�w���3���XJ߫Јѻ��j�^������ߢ����j�A��l�x/}R�l A���h����op�H�� ]�A���K�Y�Rǚ�.9�Ɇ_u�������`�|�R�K�9}-lV�1�9Xo�!S�|-/:�|b�(Ɯ4ڃwA����#�X����k5h�y�_UX�e#�v7$h����E�]`܉{�-nۭ�����s/`M+���ɽ�o����{#����b��I��s�wCb��Im,E�t=�A�o/����k�:��u�0��Sᢥ�`�,-��&R��$Qn@Cլ&Ԁ��M����l"��8`�\��_��-*���"+]��j��%qV��":쵿M����IC�0���/��Mq�����F�J�����Mx(澟ʅ?���o>\7q�������q��x��mӦy�����0�o��F��9��)�F���O�n����6�U����-#�K�ƿmvߙ!�v��7lu��Ye~��|Z�xB�T�Q9[V&�K8�� B��2�]�;ڢ�̆��w|]_���q&�6��I׮V�����(Ʋ�3�)�P�Ҏ���}�-q=l���@�N�h��'�ds���0��E.ҿ���8	}C���q���	���#O �!�qG�L��ē�Rrh���nF�ȓcKf.e���G+�Y�����Qb���>�47WNԾ���
�N��Y9�f��MA�mg����Wt��B���� "�C��w8Gu�S�jy��������7N��M'��\��� �35�4&G�6�Dc ���k���S��7*�0m�B��T�2�������I�a鶲U6���D����4Q��8y��!*K�S��2b��ɲ����Ψߠ�j�!���[��x8�\2���5�6R� (�.̀ё�aL�����L�z����Q�0���Is�qV-�%��t�Ӎ�(�+6���B`���*
@
�,-P�S��̇�ZHz��ٕ����p��1�nf��L8��� �g�hIhҼx�+ixq�b-/�G�|5�ѷ0��F��*Ъ� v�! ;���>�G7pS�Ą`ϼZ����aP�z� 2`�HK �xCulK0��_�-nK��
���f��
�Hkzn�"����$x� �.i��*��ME4�*Z���/D٬|'�w�p٬=)r�9oU��V�Pi�U���
��)�tS�����C4l��=�K�����â��rbC�/y!�툮��!o��1`��`OQ*?��7�:�@�w�K��آ�l��U�W�U<x��U���!tPr�uo���?�t<���]�<%��`p��݇>� ��@�P]���@uؠ����h�G��<���xYH�4>�2��7�Q7X�J'�vS{Nk�	l�[>�s�ș���'��X"�!I��j��<���=\15a�U�j��0�tSY��� S`�F��a'ԚEt6���!���s^�{a���⓱����U�(a��"��p� =���f�������u�+$�FzE���q]�յ�t?@MU��S��_Ң��	���f�ǐ��o2��� ��(��p��ChЭf�i��Q��+����*:$!���]�t7���ܰ�]�,���k�f�˼=,sJ(��]2���2՛>6XB�7�J�M�����ssd�ə�j�%�&�,��菶W\�4M�KݧN'TA�A��Zn�|��]:'_ye ��E@�'���Æ��󝉺_�r��'E�Kb����T����g��w:��<�����f���ͯD]�8���K�e+y"�L�.$;����P�,3�W��������g%G���E�v	�U�5�q�z�Ia�5��BO���]��3��X�̎����>m�3k�L!f8^%����� ���`��n�[`Z[�߶,���~��y|��*���`5@SP���
]:Wh��P �8Uc��ÉC�Ji�0����l�!gu~���`���7�c���K�����,أ�j��4YMo"�U�ɢ��6�*X��GL+�n�.jLk&��dF�,�)�7$��0�L�Rg=�kM�v}Ƚƿ�2��ϕ �FZH[cμ18���1؆�Z*PuՁ�*�����6��nn�:�#E���9�h��Kt����VJKV8c[�?���_�.�?�;u/w�Bc�\#�j.��7��{`e<P�vm �r=�\H��u	vSŗ'�Y��!o�Vk�h�Z,c��y�t�*~M�ZM��j�_$��ˑ�������'5�Qg����e�7�����W�\�Rd{}�NArFz5�ߛ�L��V�>�t8o$y�u�{��9��}b/�Z�t"˸���x�(߮����#�Ko���t���(K�,O��j�[$b{��H��*��kU����a:�T���(y�U�"E@|F����#,�kw�JI.1�S0��;:��Ǿў�C\;�
��&h��a1�?�_��C-Ŭ�G&��RS����0��T��]��¢Nǿ�6����� x���1�A��K�@�0���B:��/�خ|��S0�w���E:}�Kr0�2ZW�U����劜{s��:y��+Uy?�wL�����'
�?�t�VP��#ca��zx��XA���2���L8r<��z�iK�>��Q���=Wv�������l�M5|���kL���%�CcY�0�ZE�J%g��ab,P"���J��M`�c�A3�)mcb��h���*^��k���5��</�D��Z�N�wA\ &hĎL�A4�� UM��^��
���Bö	hY���&��E� ��f��ms�V��C2���7��4����f?�S��Ņ�g�t��ch���һ��H�������������\��T�W�a�钏~`R�����ҽ�ӊ�����o��ɶs �5_3��CT(D^��\��b�a+ e�� 4{�&2��~MQ��Q� ��}�v-��D�rga�z";��z��6��@L15�'}��?{h4��Z@0�UG+Ļk�oq�z0���f�����W	�R�i�|���FrnG���[;�-"��CYJ��"9ا-����foJ%g��OY���KL�[���x5�'k�����<�	���y�i%u�g-��}LCO%p&���fp[?V�[/$�}�pQ�د��fP� ���Y�ѹ|g�X�>�.�O�br�5��~�?6�$��'P�m���_q���j��:�S�R��Y��r-�;�Á���=�+���V�<N��%;�OҤ�b�2l/�o�@����ĝ���5�m)�yt��#��qv�����rP����5�
�$�*�i�j���}<�_��g'wZ&:=�l%X!9P�v���y�#�Ś�/�p}�vO���цQ�!�k�ӂ[z��ȹZ6|d��#���N˦��&�����oA�u��C���/�HAMtF��F�����~L"�y��.ٿ�W�� �kAr����:鴬8���]��LK �e�7v�<�NV�'ka�>3�
ϱ�q7��]�E���ȟL7\D^���N�G������ZG�?��X$�8Œ���=BL�xY�Ń��w�\�6�\����M�he�5
�h�����l�t�M5����i�)ɴb.d�$��4�R�k���fݕ�Od�,
� �F��v�/5P���W�6�FJ�u�� �Uw��iۺ$�.~�uī�$76��8���cQ�_�պ�|�L��&-�
 x�(��;��@wXG�B�Q(�\ˌ�x�R���ƽA��P�Ӈ;��z@��ٮ�{����{�'��X��-fK?+���K܃a��0�ު�*�a}'M
|@�F[#Oz������CM���s�|Rw�P|���� ���q O
�5��
t$�\�^sE���1�z�ԃ��2$9�`?�T����9��N���	1]�	w��A�/6��bH��M� ��%j������-P��̠�}#fϫ���=�Yˊ����h�I<��X\��� �-��Ն��VZ�5W�����)ǘ�z,[�%��C�����g*�y$����2t6��L��\�v�O����������1�"����(��v����W#��>�B�XØX A}b;+ڄ�02�ɑN󕕨� @�|�U���=���[��u�hc�܊pP���6o�1WX�.ԅ"@h�1#���-�;�EZ6e�}y�,��R"?�;�
n��c�,V:�7�q"�kƀ��-�&�98����H$�Df�~<�J�Ð�>sx�j}�o01c%t�*����g@��&	�+V�W�3^�r9�iɘ7���8eC�L�K�l����@�4�AU'���.F�vd �ȁ��C'5��XB��2T�D�i�/��g[y��$�Z�̼��֌�<T���$�(�����b!\�v�&wF����s��(H9���J���ʌ,B͊�`n����.�G�9h+tF�&����/+�23��9T�1���'Uxf=D��3���J��0ː9���e��Jp�f�^@�uxg�
o�u(�ō�ָ�.�LQ��T!�/B'[aH�D~X.�&f�Q1���i4��l��W��r�ku���.�װ_[�O@sb�Sۋ���e���6N`����LL�$�&�$��������&�3�3�e���j:	;��栺0��YX;��h#�(�mr�Y�|+f�ʌ�(Ы�B��=k2�7V�� �Y��XSB��HSo>����d�I&��r����3�.�q�k��mhקij�K�7�;�J��f�`��%�<k�(�>�)��M�+��j���9Q@�]��Z�za ��X�aA���'&�`�)n���׳��V��Ǌ��D�	��4��@��g]�� 9X��������:����.q�N懲3!��>If�� ��j���R���l��P��:TX�:�\C���:=�H���Kd�D윤��#u���A�?B8�b9�JF8��(������-�8�p�K����`�?Q�/�QCՔ�G&j���o(lpX\�O��(� �nQa��7hdMH5�8\���M�
�y� ������W7��>�����n;��P;G��Pc�eE�`�1Ӯ�����e6o�N��FB��o�)�:c����O�0���u�m�a�.��������q��g[)*��T͊��7}w����R��f���u���HA[7B�>���K�]���~�O����m���uP?<�QOOuA`�^2%� �>�B��ƳS.�AŖ��Ϡ�"`��[���?#��D(m��A�^F�s�l�Ϙ��m���q�T�!Wm�K�4�q�����9İ��Uu�[ z���H��$,�J�7w��L�}�i�K����t��m���_� ��~i'�j��I9g����Z�5�\*�C�!���
vo��������Մ�Z2:O3���O"��ƪ�t��B&k�F9�����}����m��5���F�Kױ��$��<�=����٢/��=��d�Nެ}
-�~78�����@Q߿���<���%�4�"8������X�*C��K:���N*D]��ln#����:1�EB)&C��8d�r	���3�w��q{�;��6x��RoQ�����kc2�;ǸM�V�n��x�\kv]�ͬ(kɞ�`�8������Id�]�^���D)箫�� �쨜���'|���\��MF�7�����
���d!����D�� ���_�3Gu=3uO�����Jb��o��x�V���zX���J����9�*{��৪}����[	*�D�G�CK�%`���4=�u*�id0Ow�޷HY���	w��a��?�Ћ� ��'��:%p�
��/����n��7���1�U�!��ᐩ>1�pEjy�Uy�w�iď;)�x�u��Ӷ�\Zu�۫-��O�w��d3�y��l����;u]�Ӷ����hyeKz!��JP>�hڗ-���$2E[��~C�eI3�K@R�����%%��I̽�@����b�R�ˬpu ��-spq8{�S�1�4�a� �e�sBCg�Z��e�C;�,-����b��:q@�Pџ�T�;���P���.��R5۰b��Q�*���4�7�r4;C�dP�`=��=��թ�}}B��VuTc:H�߿����1����f2�KXђX?��	o���^\�r;�n���"7�D�*}l��w�&��
�y�,� o��+\?btv	4���c�A��4�,$h�̕��$Oʚs�� ʿ�CHDѫ�"V"���4��1 �@V���|�m�`�K���LD�,�N�2��6R�^���v �Uz�8)�t��3_�Z�"��砲��jl�a<�ZC9���8��#�Y+�G�b�	���'��,�n�%c��������a(
�>M����?l���1,���	K���8�8����@�xS���j5�P��dۯX�Y�"oT�{7�@��$�I���DS�X|���%�b"�qPF�Nd{��9����-�N�Ǿ���&���/䍯<�2;�����xc1���Lw�e�p� �0^C�e�r�u�B��㑅@J� �q���}���9Q�^#8�"����}
�j��M}'M�x
����x#3BG �ņ�'�56���U�P�ƶ���!"nȑ����	�=�������7����,6�Im�Us���E��G�F�����L��iԮ���%6;���6��_�3a�zg�b�3� w�4���$�L��QO��~���"r	"�""4����X<�mt�pj��eu�ވf���Co*��I�֣@�V� Myu�Nf��B/���U�"$����:���� ��s�M�\�F�uYBek"�4؟ex�T��Jr����g�v#�f���2��B"Jq��i���F}c�U#9�Ğ܍j��A���̄`\�*�D��V��$�+��ߺ�����'���!8�>[�����[Q^H�k�HYh��~dgJ��0F����ʼ�y��<��?6�F6OXo�qǼe'��D��{���XGP����{C�ܖ#�!����W!�t�"�i�/ȱ��؎�~)���G�/+b> p�w�9��6,�	|�.x
s�&������Z��F1a��#����.5ꛠDi�&��n4���2Y:�GE����b��x�F)�6�A��Ɯ��f�\o���\�[G3�;)Jg��Ǧ�z"Mm����D����1]�Դ��,Dl��̠���>0��r�a���vO�� ���"�s�����&PrX��&"�Hs�^�nl�pش/J' ���K�e���}���hQ6~gna^�s�N�s!�WB�6k~(ӃLb5�XZ�=$z�ǽ;�[ [@ñ|��R����������(�m�)��V .8����v��9�+�z8���m�G�L|Sڂv�iA*!d>1PZ?�`�ȝ�Jq�"7��
w:I,�L}I_������9ч��L�'�ݙ}���K,p�xkI&:{@�ÿ�]�}�bc- Ѥ_L�S��G���6��|��E�I���%�7g���R�= ̮��`�F��7\�a�/&T��Q�L�pmK������'&�V�>�3n|����PtD�n�9�=��� �	7/��}H���m�vlDT��͈mE��.Zv
�/~p�_!{�t��?'�B8���!iX@V<B�H�V�<J�����:��ˁ��A�=��C�<Φ��5��s�\�$�-��l{�N+M�\��A��3��W���Q��V]�n)oBؚ[�x{C
p�iQ�!{�=��׏�s^�Ч��s0a��+���nHg�v5`N�P=���2��S�]��ﮖ��*b9t�ȕ�i+���G?5�QP؊����>M���L�J&/Dٮ�p�F���m��~����h�W���Zc�MƝ��)P`,Kɓ�}8������J���h���l�O�eqZOQ�� ����������D��_���:�v�U�ZtR�6�b���a�s�qO--�-op�B�r%�C���2'呦��ٽ����=蚤0o;��AN�
��9�>��w��[�m���H܈ղN��?rL�M;�0�X6�5C�A�;-ƳZXTĘ]F L�d���v��w�NzA�Ck*��N]H;c�(���!F��0Ǘ`�t5�{��\"3�������|���,����V��y�"��G��y)�y�L����ꤗ_ڪ"�'f�Op�,���N���}#�daU�zf�Øb
���^��^�b	�=����ə
`�e�^��k�h٣����˳��
����&y�/�Q��%{'���A��-tä�?���a����I;ɡ���N}�I�"�VtF�$ʦ� �pmW�i~�q���/��sа��y�bg�7Bc���鷏�r�O#\I �Zy�/���<n���9J�s���ۙ��(D�,�I�0R�Du�b�9{��k�"0�p|^y�폼��*u��T?Ć5u��5&���N^԰�kh���n�hҵN)Uږ���yPd]��|`w��)���*�uyPsPS�� }���E�w\%385B<�>NǬ��V�H\KCժ4�u)���ϱ��2hk�F�z�EX��8� �{�M��4�R2�c�27Xd�Heɛz��h�z�h�4�݅$��i�u2�eM�U�V?���fB�/
��>�u��߱���?��i����|_,qQ7	�4��#k	��qp�uL���d�:�E�Y���O�k�f1�<5��י���>��Q�Pmͭ�7\Ɓ�Z���*AP��8aa�7�Ѐ��i-��e"�^˓X���ϩ�-�����BL�ܕ����n4Ǻ�'�]���|���Oed�F�ߴ��]��9�d��@�r�^�_�u�-W����x��Bl]�e�o�8�XV{�4�@lv؈��Wio�O���BKMp
��</�V 0k��M�����D� ��4�Mvq���ɽ�o�M�7ss�����Ȟ�$.a��*Ð&�F�?_�&9&�o�u�t�plb���K�~��E����ᮄޏN���"}��
���=���� 
5�~y�B#�B��77�S��0Q��T����h4��B�S' �2>RmvyfH���+^c�������{��f84spL]�y�_�xhM�?}���2�U­2�Q�Ĭ�A ��L���d���E�����������plw�����J�zx��������C&�&+�����`>K��8}��E
2i=Ǉ��V��� ��P�$O�d����>��d��h ���(�>�H6r����E�Ţ��/dȊ>:�#�*�[횩��=3������Z����f�,_��Ȗ��i
<@m�w��zz�-\�u�K�I����5-��=���c�,u���& T��(o���C����N1�q	~I�ϭ��]j�63��=\�TI�
�(��C������� l;4�i���)C�k}}CVrj]��x��G����G2?zFS	�[.c������Ep�M���+*�崸F:H-���6(
K�*�|kz���\Y:�6. ��rO6��j��^Xbd��^B�1@�����u�86�%��$�ո�����{�``|��0��1>�a���w0�:/%=��ha��Z��g>����p,{�������r��O=�jN�Vze���Yw&ɭ�%϶��[�<A��� �n@��4�O��Fh�*���qo�D��� �(���mB�7�j��%Eި	u�7!Uj��Y.��i�좂
m�x�r��W��~�Y�4�<�<۲�m%�h�k�%l 5l!��s̕�/[�
�܉8w>3Me{vHޓ��O69ȫ��k�:�Juj�����Ϋ3���ͬ{�v�#B��Q_���w98Q�۩�)>=�%ro4��BFOE�V.z3O�`Y{v9!<�}�޾��o�"��F�v�C����eXJ���z��uU��-��cL,rf�w.��0m�K �쇉<a����_XM<x=�6����A!sD��~a�FА'�%�`�r��6����o��!;���YE�w=/lOT���ApZ8]��k����	��ܽ�*�9C��ӱ�,��FQ��F�y��a��*��մE���	�����M)���`����Whȓ�&Ez{
��A?�����7y!���M�G��%�d�[���!^�΅��R3�)e�iZ���ЉiC�i'i�}Z��*�v�6�6c����e���pX��`�ʻx}�dc�t�j�x�Ƅm���/�������є��(bT��~�O�"$V��3l��!��Bj7��1������kqu?x����=��Χj�8%/�=�ߗQ�Zz=F�&QJ;rh6�Z���~o�j�z��vtV�^�ڋ(���X��+���#W��s����6��������(� ��~)A�v�\=wB̗��;@"�"TL6^S���ڥB���	^����y�Ǽ�}gj�ĀF ���V+\�����0���,}96�/.��D��O�:j��LBk"�a��x}w�w�lڦ�4�p����?���H�����wj\��or7�ĭ?] ���U�&vA�#���329�x%�}��Xg�i�����O7��I�Q�<�]�<�e�~���D� ���`7���2"������/)���B��Cb�\g�PG�?
���lPc��h��-�U&�ݎi�%N�}��|꣦����}4%�����`���+�m�]����8�u��h_17�p=��R;V��p�������N�Up2�X/V�>��ey��h������W�6� ���"�i������������dRoqj"���]��8`ٜ�+@ �Q.��uW��Y�d�A!�b Nݭa�lM�[���D�F��R��bp�!����" ��F#�k?CZ�T���z'))�=�q�07����M�V�Ai��$E@5�B�Xyٓ0sVl}MA��F:'�ʡ8�_o�Ӧ"�8�v��<������6t��9�۶L�_�1ɧT�mjr� \T�.��������վ	����o_��6G��W��ǁ�>
FBm��r��Hxo��yy�{��'(����,b,�n�N7Dc�0�aa���u
�՞�����x���{��<_���K7k ⼒B�Fm]����'ɖa���i���ѫњE,��З
e�
�6�����BP��OH����3����	������X�U!�l�p��%?�P��x�`�����f��@l��.�6�8m���*5�}���hT� Z@n�U��n%��D˸��Oy�]/C��o~�}u��/n��fҎ�9$�#���%�Qq�Wh��O����cX�p���@ތ.<�T
�hQ�pj��]ҠI<F�d6���)(ϏԮp��t}�x��&?#�x2y��m�J�J,��&Uc�����H__DL}�SQV8d����:!ٳ"o���Qn���|����9Y0�2�`��}[��F�9�)�&6~]��{y����ܷ!�A^���4���=��%Q{�j$�7\6�Z��� �Z*�<�e�М$ښ�%G��S�+I~�t\�p̼��<��Um%'��eٸ�vtbo.�_���:�
v�����1����)�V{y��!.�?����3�;hú䃉�]��AQ�ը3���w0-�a��=�ؒ�øc�����C�����Y�Ȱ�ك<p3�Ӯ�"�:��;���Ʈ^f6��a�cUJ�+��ޤ^�v4�,�A��,Oys�DEc��"Y��1�O�#��bN�I
m2u���9 8"�K�P?&�H��b�C�/�wk����CtP� ��Ӹ
@x����R�o�m�����%9@pK�^N�p�ǡ@'w��_�������U���Ԕ�L��q���x]��,Za��v�C>�$���P�
0�*Wpy~�������:�3�1	N�n +�����<_��}� Оռ��I��������X�k���8��}���T�s#4++�)�V�Wkb7L���.I)Fq!ܥ�t��'����N��(p�o<5�5�b4�S;�ը�t��]�22�-��p��Kv�$(�����̞G�}wP���)��Yz )cq�;J~ŒȪ¶�G|Ca\|�pU�p ���gL�Y��i�R���z�8Ҟ����Zj�e(x��߹1o�q�?.�������m��[���#��"��i)��˃�I�0u�;2{�n��(bKT��"9+�eb5{Z�_W�C�%,/Wԏ9^�p���=�[ן���鵢=1h���Wü�	�s�X��,\-%�k�)P�8y�3Ѧ8�H��2�0�'h���'>��ng�dӧ��\�:���6��8����K3��IjUXT��?w���콚Y6 ��l�����A�~�@��n�z|t� �[��w� ����o�6Z^0��KS{�$�H1��jr�e�gr�0�WSR��T�&��X�k����x�y#�m�:/�b&�R7k�IFi��i���
j�x�$3�Hk?�pP~;�{ٛsD�G��mn�)���q~7m+=PxLj$��)y+%��w�sK���}&B��_�DM"^���t��X��djT���q�����٣kh��yZ��j��]�iW�j��U2���٫xTń�]`V�6"��{����ͼEL%�X��|�Z>3sX���6xr�GTմ_vF�m�x�-Ӎˁ* o��2���t���0�����GhZT�9��3�M�e:��tU�VK�([�9�t��l�q�&�{�s�=���d��)�Y���s��YAٳ�/�|�X�Qp%ET�tA"0�*�I��j���߇�CdUԦj��v�����%�.Z�EV"̿�9���e%��=z[�3��v2 O�I=���#Sb	��w�23�`��6W��X�q��PA4�4�׾���x��]�P�&K�;���j��b����˒��L���^�c��Tț��r��d~�k(�i%�y'(�zC|�8���Yr�n�9����(z�PA�]-��sn��J����:~�Aݑ����G��������ps43���$[�5�P��� ��&��&S���fu&�S$GT��j�^\I������~: ڎ�f���q�d��SWՏ�F�1������a!��^+���a5��+����2?X`/9H�Շ��Z�nȶ�2��ax��˪Һ�ş�+J�M��L�"�,�꾮��&I����5�õf��Ƅ=�̘ q�a�)�3F�s�.��9��]�q�}Esgף	:��]�L�ZDp�Zit�qrI�;��"x����I�.#!��A������l��D�����ሩ���A^�X$]fL;�9O9��'�sۈJS�ݚ��h$���N�Q��+i�[b�t�2"~Ζ�@͛.�]n�~�x��#�Q]{ +Ʀ��0݇���h?�8&[��y9r���?H���Z�\6桰c������j�4g�?�O�ST�u���e'���S]F�ko���+��5L�Ѓ��-��k{�����}���*x�8�>�����̸S���U~&���7v7w��` Uji�=�+�r��t��wp0�p�����d�
�V�v�Gi�d�?v���������|�e&��B���n�'���k���~U����[b��LX�>&ˆ}d��~� ���g��k�����0�y���7ݜê^o}ż��Y�ń@s%���,�'��3�e�0�4��������5�0y� 8�Q���DԀ��:g�;s��\�L�a�E�0�Hfs�b`�8��Ɂb"��둄�x�u�Cv��2��Uⷨ3IW��a�)���*��f���t�}sI:�*��4�I���"<�6'sx�L�\`�K�p�	���[��B�De��F�v�U�| �1����4���#��0�|`BZ[u�E���SkKL�5���Yǹ�T�Ӟ61����FLn���%'T���΀eG�+_ř. ���ֺ
���/lE��H�N�� ^�q���k�eύ�K���;_`�S}`�	��p�����0Q)w��0���^'��N��,O�gUW��3�բ�G[!���q�DaKy�xk^�9��a�q�yV#�l~��چ�G��������{�J>g\�tk�ְ�ua?/��xB�[�T6OV������B��<�_y~�>K�bTk�U�c��)5�,�99�Ѕ49m�z�P$x���f�U��e3��	7n5���{�U��������qYj�4Ҽho��	���(�|8�<��rA���:����z$Υ+{,��d��	�+�WjhƔN?=��Jo��� �@�H�e���/�^����d��h�H���Eeo���|�x4d�Nl�І��Z���ȗ{h����w#��>?P�zs�<kk���� ����C����{T��C�*�Jc?�*D�s���"�HtxV�6��x�^�\�=����Xe��,� ��U�=Xq��u��-=����%�y�O�t�C5�!!F��CV��E��o��V���}�����zg̎�
Ȝ:d��0��԰��gT7f�~$������$�>z.G�q�O=�2O�ގ`i�E�c�u4P�~�!+�
�ZD���i��@3`�w]/#4wd�W�{�N���&z���s���kb|	�~i�^�N��J�;�����K��G������JJ��{�rΖ�R6I�^W�iD1�XV����$���Z��wb���G��us�2��I�/���l@�Kbv�@ݕqq�˗��~�ç��qk��2��m7Ov�Na���B�z �Sx�`A�<Р�I6,$�R r��I�-GŰ�:J��9����]�djN�ќ5b��J�ɦ��,&�p�~
[���d];�����5#?���%J�o��m.21����X���|����ݸ�4�rTS��
G�<TTKg�0)�J��������<8מY'�$��T|��t����_�jD�"��� �_��X�t�L}�Xc�k#$9gX���6��YPF��fz��O�ۡ��	y(��@��D���4v[%�)k8d�-);���au��_���5��.�sMFY�y(�M�Q?���xm��DT~����x�՟@�=>\�Xx=ޤҶ$��]�'p;�z���-o7��&��8����oks<�2��y2��i���oTM���q6���̒vP3�%}�-�j�Gj�*UR�(,�KU�B��,���p��Q����E�'wC�#���	�(V�*c[�x���04=$�\84WƇ��/�xŨ�DHQ�R@����Q{���җy�(2Yچqڝ�+x��ũ#$a��D�FϘR@ev��{�P�6,>�ҡA|��1җGx/��lI�Cf�FmG��EQW�J�f��j���kt�%����;~�@����^)dDt+Y]����mza[c7�pʹ�S5�1���n���>����s;��3�����R'&�p�7ѱ� &���Is���)��D�@|{  ��`v��i{gYb<�����3l 3k�Pw>��Ke��0����Jİ���Lnee���8� �I��a�C�/\��#�x\�
�Nc2� oʬ����f��Ktۈ�Զ /�u#����8l	k�q�X��d;=�4�ie(�I\K~
/�-DQRx�9i��b��Vj��\�+� �q��n��FV j���f׿X�+��&�������D��Dl(��Ϟ��#�uٖlky�� ����6#AW����u�j�*_b�x�.�w7���m����Ĝr���Vԭ���u�X�U��5��v�$�f.ǻy�{��a6�oҋ��qb-��4�H+�x./f�NCy�I�{q�����;���>�����=4K{�1u7O8�����Ƿ��4���-�@�F"����{�.�����}����q�ݪ��7l��m�r�`j����d��5>�!�'���'!��J���ۗﮥ#q�/8,e�ܡ3��5(�cA�LG�8{zMɜ�X:*�^kD���)*CEn�d27���(�`v`t
��9��͎��s�4h���@�'����Q�	 6{���@�8.�<���G��3%\��}���������J�����������Y��t���&��^ج�����܈5L��ũ�(��-��i�b������bt� /Ͱ�c��e �]} �.�_�0��B5c2܀�3��)n�{�[/g=*u��8m���ZZ���§}*�ΛcX�h�Ʊ������JB�w�����@8'�̈*uU�����g���)F���9����7�x6#��j�S�>�d]�8�Sps`;)OSZ�t�*`=�rXɘ��Y2�wlHʝnM���x:<A���t_�}�;��3;��ՙ�(Q�M��yL9��sxifj<6z%�j9AeךA��?&3h������(� &��H 8�r�V|��I���]L�΋:X��7���7���zF�^k�����WL����GǬ,kr���V�sTV��	8ٲ0��o-�8HX���'����� �"T�"��Z�Ú%�]�/�^�SK��� �@8D�/�t�M�ѧU77����b�O���]|�SC���Ym�*���rqQ2���&���K�
6|���x��� H`CR�"�:J�~��C�<0�Ej,j��8>%YO��i{�$E�P.�?��MEӼ�\�����Z߉�<'C;U/��i~B(J����6�p�lg�����v���+CE�^�Ί(,��~L/3%엪����/B���Ꭹ�U,;�����!�~���z-����*4�T��}V2cg�"�%_�و,����@d;�)�H��X�Z5�`�6y�X�i�ᐖV�rX��!�W{�+��r�1Y"�J'l�˗��?zx��P���fj�7m��p��v�#Cg���u���=�lM�wv�&�>ڀ9H��g*J��)bTg�"#0�� ḅoT!z'�W�̰�6�����H��/Ҵ3�셌R�9�\�J�,ڙ�K�>��!�9�<v#�@1����پ�&yJ�vD������W�кs�����$4.��Oڋ �6��ۼi���|XC݇�jo�POD�p������񘠦Ƅ˱Q�er4��)v �#�.#�aʕ��uT�ii?��.�匮��A9x�P��r���Os����Y�~��� j�_2H}���o}��Kn�W��%���ρYsfG'�я��ىC��IC�k�R�`�^ӎ
?�7�t�0B�b�*w���A��\���1ۧY4���ƒP\�%�zMe]�d|��h���v-UR�zj��[hY�Icqf>.�Z��X�"4�#:���i`wh������]�`�>�QL[�,�%��|����͑��P8E�Td�|�U��I� ��Y�����Q~�v��IT��=��;�Õ��`�S�����+�K}�e�a��n�f��܂�}�I� �}H�>CZ�k��wG�3�#THI��S�R����4�#��NE����d$�����A���5�Ւ1�@���Uĵ����Ĕf@�K�^�����-�Z���޿�9ƌ�FLv��Jh}�n�Q��oI���s���&[���u���`t���J[
� 1�*�O儢�^�`�����g��_yeW����L	�������TS*�eN8iZ�q�N�д�T��١��f�v��U�P���N ��]�8�&�O���=�q��տ Y�s��{+"�Y�0$�F�CmĜ$M�G �k5�P:��-Q���Q�^���*�C��y��)CVl2GٜV�;HM�̡�#/:2��T��ʽU�<=�h��yu+٤A�O���p�{��Hoj,�w�zk�\��/M�}+'��r����}]�� �?xu�Sf���Y���F����#��
_��pF8���>0T>�\P���$��׸!�6�5z��oI���[�f��L\���k'#�$�E'IG�}����qj�Ÿ�<�lKtm���t�VX�L#�u���iM��,�6��4]e�lh�[^�b�[�����*	�����L ���!�oE��&J�s*i�!�����]ġ�o��䡇��Q�U6���q�?4�Jp"��0ݴ��;�� ��#.E�|��D�$�
d��j�zM��_)�������jk��E�`K84�;;9_�2���}4g����LLAHv��U�blߣP0O�����1���9��Q}�D�K~[���M��3!򚯩3��h��]��j��q�$�Yݍ}�ㅨ�=���4_Χ��u�>��F$A:��u� ���0����x	p�Q
rvk��R�v��~j��zU�I��w�~-�{j?�Z{oҿj|�Vj׹��w
Y4�7��BV�� �i�^:l�VF:�Wy��j�Ӧ��M�y`ਸ਼/�^��&�06b��Rix�
��,<��ɼJ�
�q���o����c�_
�F����K�h�s�Żާt��v�#����Bam���ӶM\��¡�ߍ`E��=J';A� }�%.T�˾���Ӻ�ja5�Ͳ��|6��͂x8���E��f�v^3_���G��u�JI&8�A�C� Q�ww�b�O�YL��W52��8:�&��=�2u�=�#�zg�����6~]"ԡ�1�u�<�<Ύy�Χ�]� GK@!�X��͐�{��>a{���8/�\�pG���F}(�KԻ��lp�0J�&�_C�;j����l���(s�Um���-H��F$[S� �6����_���G@�������4���>;�x`y�����N �D���ͽ��5܆%7#����+J��P���E������֮V�]�/YI�E����w,GƤ3�h��~sְ�7��P�E��4)��#?�o����̨��G�O�߫(�Vd����$���f۽
���D�/��7����e�"r����7��HV�&i:����sp�,��(�m��k=UET;Tez����a���`"^��an�^݉b�L;YC�6@L���N6S��}|ⁿn����*t�A��P7�Զr<|XU�	����U�D�����g��ɦ�d�!k8i�L��E}�Y^���]��,iIs�n��8�^|_�?�'w`-:+��!5��ݖhҜ�)�bK����F�G��;m�O�v���p����`��M҂?*�#�nfA�;��g+n��t����g��xd�)��$_�<w1! �������s5�ijc�o�U�V�����$����t���ę{���A��e�Z�����2�H��W.L��W�+��2p�@�
	1�ܯx�t�4F�If�,�dc���H��a��`-%ӧ �t�_
����4Zq9�b �ꗴ����������lv3���sТo�kldp�����O�M?3#�b�ۼ?O�
XDd����VI�q[cDײ���s��١,޻�u[�* ��Ѭ����=��0�F �u^ e����|
\NTc��_���ѧ�x�X3Ū&I���7��R��mS��;���Crc�h�v��yD�����ΉK�i�
�!�t��������~)�-��]G��Z�i3� Ͳ����:�+�$��I�hv^*���]R\�"�!@o< ����ڛ�A�1a�"��7\W��0g�;�DHo9��'囙�QX�s⦋øDy/��-|Vp"C��',Wx�����c=8��`�'��&F�!o�XP�9 �^�,	GB����ܨ՚Lk^0�/��t�=T,ϲ�w��z�3`aDےq�Mns�~����l�8��{�����;��am�z u����Jf��;���`*4Cཅk?-BG���a�i\Ϫ��xG�7D�v[�#*���wb�'{V�#����1���~��Y5@�"�A���̆f�pV�u�s��>��}�\��=��QX|P���vV��6�97h�s����1a[T9�fv +'���`��?��ឦ��\eC��P�]��:[�}�~Ԩ��l��\�)b�h�GR�kY.�8�q�2/������LD���SK�Hq��Ǟ�{��2O��䊏�V�,Ejc���5,Z��#t�mQg�~#_nV����/kYX��2}:�S�-͆��n�c���˳s�2�PBnfA��?�\:������,��� ��0��LX}�y�晄Gn9�g^����U���t7K�'qQ��YM���T��:�uv%�B`5�Ǻ���V6x=�hK[}Fі	�x��@�|�S_���N�ra��O�tD��m�#UN�3���.��G�p�x�W�)@4�x�QZ�팚���)c������7�ߊn��r�hv�$�\f�����ߊ����F���T�٘-Ӗ�ή��v����V�!?��Փ+,��
�C#W�=�������Y��L�Г�T^r���m�� �>��v������E�8.�S�q�Fj���~��鰞���a
���.cv�&!b58�n~�ug�/���$N��4�"k�T]�0E�W���ke6l-}+���) �;��H&G��+��O��r%��2�z^\��+M��T�9��n��o���q/�{�T�v�������W8#��=�W�k��JD�n����k���M(;F{��s���A�!vyϸ_�?�N��>i~U|��vE�� u�b��xߞQB ��C��qj��ݜ^ik׻HM�!Xv)_��,.���Ƿ��V�lqž85)8�Lu�zބ�B�5jWc,$�fm��j�1��!�*����
^�'+���+G۱{<�$�j*�Q%��y5<��zO-��Q�ʓ2��R���B�B�oC�5X�yjAy1_�Z��Ӻ�����;	�-u1+��k��[e�n�]mj�d9����I����i���?B�n<��.�8 ��t���9S2n�3 �?��clK�3��<.5�Ip��A( �6 F(��
���L�R�N<F����}��ؘ��ԣ:�802b�]J>����p��E��{D&�YA�VrҬ/��D�C	���ܐ�9`��w�53_�
�����9֕;�N�U����W"�\�1���GQ����;&�(��2�_	&���&� �?��z�d�M��If� ��9Yϥ@nI	S}�ξ����w��S��%M�}?��L��Mc�P���,J^[0l�"md�Y���gV�p
�MtTz[n����4�bM��T)hVQ��U�߿����Y(�fp���U c��"�Ǻ�Ӟ��<-���_�,q�;��1r�$]�]�Zd$ٴ�ƫ�0�j�͵ȥ��� �W���RJ"��(]�fn{y�	Nޜ1���l��4-l�e�54�����-���l��_u���2�'L����1�S`�C��!�1����2�'�U�S9��y�����Z��&��m���w�-g��H��|�����9�f@���F�-M�l/�UH
���;5��L�vb2�!#8s�	��7��;�S��#o_Qx�1J�J�y	�;��L%��y�������!��˳�`�}B�����pB���8܊s/�- 
�
�B�FH^Ǭ�qۈM�W�2���R*���{ȼ>�UR�X��G����7��Y
����]i<��?���;�gt���s}Uٱ�U���)R�V{3����l
��U���K�p���Ԭ1��s��,��L�l���2� Pr<�&����K��������bJ��v������p�Ϝ�����&��:M�d�Pj��B�FD�Lm�����SzcK��D!�b�?�v�4y]x�4F��yUɎ�}�񅇫�vVP�����5�G�������������q,'���Q!�;1s�Q���v�j��6E�=���Y]�<���ۺ�RX 넗�ʝ��GUY1�AJW��<����R<ixS��=v4Y�!��t�iW��Q9]�,eQ�zg�c�����x���e|�\�����P��3�ej:��m�F�����e��\íS$�˨�N���чD8�V� &N�����r�EI����.���>T8V̠�LX_���{����AxV�����zs'��nB��!�-Z=7��eF|af.&Oz@�A�]1�����3u^������}���ԃ�(���m��
��Zf*�s��*|������1�9L#8��"M���=E�5/�K¼G'�J�dw�9�Q^�.A��xS�+��(�� �]�[8-)pz�o�o9���X��{"�ZG�ܻ;�n-�&�OTf*�ݥ��[�!.M�dLN����@V����bn��P*.���Ʌ~�T��(}��� #�X6�܎���E�@/��!�܇"���ɱ�d����극d}2 �¿�N�u
�ÿ�->�Ğ��`��!i��s���`�:s�4���̘CV�S��E�7˼��E�p��ke(�2W�$0ڮ��*����'�6�?�uD���D���l�P��T]�84�]�V}���<Qq��C�?���Z��i_� ؉����ecn��c��Ro��iy�I�;�D=��8�~�ny\��(����`��[Қ��bL�>u�����_=&��b)'p2��r��������Kq�fU=��ޗ�F�ˀ��o��=gl�4��1� ��ˀ�x`�ce�8�w<���lI�1{�����n��W<әѲ�o&�J�^��)�Ojxj/oT�s��k�moѷ�0�`���"ہDvM�N�}Q8к����>�0%��'�w9!����#���&����N���:79{J�"����B�V����M�����T�2�t�oa����K�6;Q�<0{�J2"Kp��'�J�M�֔�9#�~b��'�}~f
@�x�� ���!���N��Z^/T�64f��{w�?� �*ܾ����+U�l�ɠA�VB%3�l�J����m��>��"V�Y��v4��yȔ!�e�L�e
��>��%�#�I#u	�t Z�;2�R��e��_U����H�5u�ۚڪ����B+��4Uo��CV�;ւn 7�X���\�]|j�)p؜L��a�%�l:��ڔ;C�,
~�kW���j��`uV�BݤU/���8I�>�\K��hE����!����d����c�1�/�n�oHX�vW���D��m����4�uaW�sG��:����-�q	D`ܙ۽��ƲߏJ�7�5���s�LC�M�'��j������i�Ze�v6�.<xCg�2U���H$�2s��%��Y����'Z�7��f�'7��Y3!H1�A�0oݟ���f��dʓ�U��=�o��>+���UѵUC��_\��X�9��[��AΥ(�l�'GCř.��e����}o��j2a��~�lɠ�*"�v<��IR���z��"�g�%��BL/ldb����8�S]߀��(c�|�F�L�O$G�;�5u��|����|�z�;R� ��V�x�K*6��-�q��c-ؖ{, N���r�:�K��~ �S����N{����jTb�&W-��T���k�����EN�p�k�;qOt���j�ԮN����'�ٛ%�U7;9�PDP�zۀ��++~���D؞B�}��Ԅ�&{��g�[�@n��Tjٵ~(~j �˟�_�?�e���@B����l297~Ĵ����>� .��mG����ye�n�g��ݚX[]�d]��¡�ˬ��H�֨���e�SmC۽ye}CR�񡳚��$)r8�qg�WX��P#JN�PoޑT_	�:�Sc�ש����6��
��!$O�XKO!�����%Q2���9i��,Pr�W��CYZ��~A��R ;l�
�xh2� %�ބ:tVڷ&98�x�Z�]{>��!��ѿ�h��	���b�q&��!ċ%́m������w�����T�r�^�#�o���5�X��8,X�%^xՂӻ��������q��4<X �j��Ԡ|5���Ԍ!��b���L�:��h!��j}	O��̔�':�9g[�o��r��p�G��&�	�`dQ G��}%B�]\��]�Jx��;������*gQ�e���M�Ö+��H~2}}p�;�[�>�m|%��W˔Z#8pH_M�_�� �c߆Ch�'�
���tt��@�Vo\'����Z��S~�ܘe��3�Lz�_��?��B������,�(��Jfc5�`���j���@��<3�v
:a�+>�C�֡�)����05�a>�|.�O!|��g���y(��A���;��:G�0�[-�2o#�z�`}SO�%�̄P��.�ž�\���6h�-bf�����g:�=�#�o+s����0����8Ḅjl$���^S�I�:zA3����2zV`7)5�DD	�
������t���H�s�.С�{^ #�0#b��2O?��
5O����Uh2 �$:W�e8^W�Z�Q� !#fg�L���}-���
����� f�e?b�PU��
���E���~c[Yu�~����+�|��3�ȡ��,�q��+���鑇�8��L�?����!^id�Q��߀�!m ��s�d>q�Iȭ����œ�qK�[Jb�Y��Y��S��"�U�;������Ó�Z�z�J0��$k/��L����" .��\WR-[(�����*qolHwE���S��u�肟�C h�A�ډ�i?�ov����:��cP��B���3&����J�Ϸ"�sH�5���lឌF��|G�ͩp/{ٵ��-Pҁ��Q�T��'�+�ߕ�S&lhS�� ~�j���8r&��`�@�h�������K��5��L�G++jTj��Z��R	O�G9���ޫ|���M;k�W�Gp�ٸ"%���V�^{��W-��E
[�\�!p���U��3��F���)�U�"�����i� ����ޫ��~mL=bMHL_�E�u�XvC	�r�[�`�L��ϡ�y���i�+�@I�;;Wrf�!H`#��7�Z�eW��~�R`j��]�_�??\z^@��@aV)`�hd�r<� !Z�HXg�H�8y��xe ���O�q��F�\�՜��Ż��_]r��vˢ��Jh��_�j����[�벶6fObr&�K�o޴0|���X[���+$
��I���i��5���:	�y62�^�4�E�l��,x�H�ġ�9���wHC�v��U*7�l��f�QP9��YtG�S����02�kA�
��Q���_��9� ���!���y��P���x"ex�@�ۣ>���yكC�D�X1�8�\^����Ѧ4
��o�u�Gs�d���̕fM���gBN��`��`�{e�*5�l_��c�**>�W�)r�v��Ey����;Mr�v��ВA���.��~���O���{+�1��I���5�Ԃ{�/˰S��E7ƞ���#���=uPe.kϨ5��&(�7�zK���ﮍ."��s�$����9�e"��A�[X��L���A�`����9um8��/���"�����O��i�,i�7�w'�=7�^Ⱦ�S7�<	�p��s �ۻ`%y7�r�򕨿[J��FĖ�0��w�M�-�x���I�OLՎ]�~�ɂ�E�OO�)?L��5u���)�2���XX��Q&��"�&�A��.� �D�v�䆤A��@!z 5g��e*"��9��?�E��P(ԅ��b�x��%��^�-P�Թfo�[�Hmp.�	!d�w=`��`�mX�u��F����-������g�f~&�hH ����+E���mH�:�Y��ކItO��+X|��H��-�:ٵ�Y$�o�Z�-���Gl�QU��*Ր�jE�����.��d�s�-�9s+���.-�1�
�p�t�-�Z�k��� :���m-~s�g��$;22�`x��D7F7Lю���(n�����6?�)�ּ�N>���I[f��/h'gѮ�"��%��C�8�+P`P�`1��嫆aɦȺ>����[h�U���J.;���H����5���})M��w'�[�ܛ��O��[��ϼq��E<)(�L��oG-�� }ї5�72y���Aß_�T*u�*E����w"G�p��Wo��Um>?)?k�b��.��,�e=5�k��(�O���-�	[��^-���o�r����г��/���J0�QU�_H�Ǉ@/�0��������q��P��Y�(
��qq�Z�]����@�A����� h��@�z1�� �0KS�1�i3��|�g�q�����{�I.��(�R�XA�ټm��g=eF���vv�Y;��n�>
�΍��5�U�k_���?�ꢱ�ݏ��\���D��?��h��`�@�a� )eꥠїA��n5��'xރ<�
Ĺ�]��p���8ks��х���P�WC(�Bڤ����@M��/�dwXQ�fF#��f1]�k�kZR����B��O[��Ú�8��Z�1Φ��E��F�m����W�E
����7R^�v�ZG���goV�LJ^Í�m�R+P���ۧ�6'Y{Nң�Eb�v�&+���k@xĄ���	cC��"�9
�!}2�-xGDܼ1X3y����>��b([\�%���~e#���=*�y���fcTe\�M��[h!�j���i���bbpbw��V�<�ѱ�'ʹga���/�A����l�ėF.��������p	V����r7]3Mȵj�K����Wm?,��	�.7�sqm�^:o��<;2�瀱��UW��c�9�ݐ�Gݏ��Ш΄8bL��u������R(.T<�l�P=m%�$��c��}5�h��%�ƻ���`A	H`1�죑�:��m!7�X�
; A��NF('����;m#��r�ʞ~Z�=����̈�TA��ג:&H0'F���^�!�\V��5���sm�k�tax���1���l_��0Ų�����R`�'����""��$���:K�cD4ٹ�E��~6"�6��6{Hܜt�)r&X����/�+4��g_ʍ	ǻ=z�0�K��
�A�?��Y{���	��˟��Y��-{��#{>D�@nip9�W.�#n�?��ʹ|́�uo���m��6�(D��q���{BL�� �w�k\fߺ�z�EA��Sf�M��UaK0�j�%%��}I�<���n�E4u���Y�@2� 툆:�yGſ_P��]��P�
,^qג�뛈����4�p�ش������l�b��D��_a|��o��h"��e��	����Dl�Al��u_��>Oė��18C�Ρ��4�.�E� T�ME!H�Bkk�a���u}E)l3��q4��P���d9ڊ��nH���f�ӈ2(/�Ά�%��;p� ��gI�mS�U2��DU�q��ʥ^Qcj*�2�%� !����l���G�����xQ���&����~*�uY]#Ժ�ӕ_���k͔y��~�{����Th�mxa�q%�M7�������c�p��J=˄������>5���d�!�8����5�Bȏ�8k�bnV�+'v�Pf�v�^r$&C�/�v�$p���j���߰�����"/1aZ97Eb�+xl6�+���(��JZ+2瑨�k;�g�"�l���%H	*Mc���k�ېg�//i���=���ö/���W�ɤ�a�1gT *�=�p0����5(ɑ^�?���u~��%95�X�82���#z�.mQm=�ub E#k�1-�y��;���� �N��XZ�[��j�N�l��
������hn�j�"	���t�������r�;ؘ�"YS�AM<�%g*�Wٿ�f�mg]�ED�e��"�F�j�;yH]_7�P��C�����@���@�	�F����|�1�v�|�u�W%�ķЉOv��0RG�T��ʸΩ(,��K����{R����
I��?��/&�s���*'J���({;����3Y����-��L�����[�N� �:���'��{[Izr�'���vv�Ek^wx������RgbVel�� �Žb	���%�4c��쮼R�h�.��m�7ϓT7a�I�P����*�:�
H��˔�"�u�D[�~�9R�Q���(h� .0��ɽ�ng�
�ti�ڞ&��R�+�k�}&��3�L��b���Ҝ47��T��f���?v��)��ӽ���g��Y^��* �\�c��9	ۍH�>�?�m�+�����Q��n��MEǮ�!Ά�����7s�s� \0N��<��_{v����]��L�B�4�G[�-8������_�`��ԝA�ڨ��M��\�����R��,C�/&%ӧ�g�^�|g"�n�Ǘ<=�E�%��=y,��(�jF9��Y����kݪMJ�"��L��.W���N�^���ā��,K����Q�������e~�Iy�Umoz�_݉�>�l����Ʃ��RS��(L
�o�>�:���ȁ�Yq�ı5g�7e~���G���d�B�&2�Q�S����ݔ�%@N�,Bwn�%�M�C���5��c�K��R����v���nʷ��GH��s��}Y��Z����;��5q�y���_NH�e����q���彗���E�8\fG1#� i���$0t!~W��0��EuN�x)�(���zN�5������[�	#���͟�+ܽ��|���}0���ʟP���<���,�\	0�`�#�ه����L��������Ұ�Gzr��=J�EIqJ_\t�.�ˎ
�pu�Π�1��6�`���j� c���X����y����A|�ٝ��􂔉���ΰ^l��5�&9�">�L��j��l�N3��}��;�zf:�·(i����ݡ:D��²p��k��q���/��FBϓ�NN�y&i�@� ?ޤ��Y�pcg�3O�N_�8-���H�LѠo�Xх&�2U���-~M?VX?�ѽ��HlK�ѿ��#_�v�S�vŌL/����'�����b��}�d�݁,��������Ȇn�/��&�����{��3(������u4 UG���+d���``� �|���?߉-��h:њ�+y`ߜ'��T4�M��4f�+�o�V<���x�x�LQwo��2T�{���%��۝��E�Z���2U M�Mȋ?l���=�[�~�L"����x6;lVu�Fa�:��{w�˾��a��2$ZaH�	Zi��%,�V��T��0��Y������C�p �r,��z��o	����h�p�"��:]iF~/��D�.��R�ڌ�I�Ca�#���k���I>�оA�8?��Z�
-ѠW��U���^�7c6s,�4]q>��o�ZE���������������T���p�"��i��0�f<U��-��6��a!�g��|�5��`{$��x�P�!��6[��.X�&��4}w�Z|��нs=�~+�����;i�=qy+�W0���EuLLU�&;��t��a�<�/�ǳ[��s�F�Q�UpsA"I	��+�Q��;��*�v0qي����Yۆ����m��5�K�iy@�%ļ�-&�F۔n�أN��+Sf���	��'�`.|�*�l��*�Ȟm�!��A���HC��c���#"~3�VjV�7�+�v�f�=l������[.�Dc�nom�A�z�Pn��[0��ñm^F���Niչ���Q'�6˃X���@��5ج�T��<II�.Rv��Z�K��7O�Z�Ro���J��<����p&�(P�Mdm#��jQ�����Wu�\��<.�׭$����:<pGW3q��M��r���:2e��h��e��w��:D�\�D���Gn~��d'8� h�z
\�H��ZUfzr��\,��F�
g'[j�<���:��8w��t[���ژH��ȈQ� ��BS����Q/o(��h7�cS���rA�{׬g�<�����~��0�ȿ� ���7�к��w\-�ޯ�S��]!뇺���܇�VoJH�����-5B{v/�|��b���8�����p��h���0�Tss����i���"�d�ؽ��-���*&S������=�6t[q\��?��.H��[�V�
�>j�B���)I���G�A�X�%עa������F9���4�;�L"`��ࢬ�E
��۟���l2�K� �I��k��{֕F`b!(�5�.+�i�CS?N�������~�>gD��$�ی�A+�d*���f��-�{��W`[�e���v���=�y��u։��tW`��O�D�'p�������
�O�ڠO�V5�r�Z2+�461����#
�f8�Z���P��h# Eڊ�ܼ/-WEuJÑ������(̄փ�'�(w+�;�i�/�3uz�%���r�2�^"*7��ص�Czĥ���6{�)�f|�n� (�b'�������,��ۏ�
�B�F+R���o�m��{�5�'F�;�;��g�0X=ш�l#�q<�o�u��e�I0FEH
�X��!�&�W3�`��>K��
P�S�M�,���!�rR?Y�u棎�i��N��w*QM����i����:_m��u��~��ozϘ8x�4Z�FK��L:�E�e���B���Vp�����O��}��t/��� dP�G?*�"3TV8g��H�t�I�{�E*��s�I��0�V\Έ���I=�~1s��(\�o%,X��rp��W0���V�Ę|#��b6����_�~{E?���lW,�Q�ǏCS����(��ܬ��jI�M�$#����;�&���s�H��G&eOe>�	��"��o�z�Il�N@;�fN�=��_R�W�r�����_���� �dm�K7,����-H�,|�N�6'ٹ�����B���VY�'(g'�v��f�BP��"���6M�cc��=�<�}� �HL)*^
U��p����G�h:�b	8��l�g���M�x�+WF�+�0�}��`u���c�>�c������Vzx�n�K������NoO��`?�8I��BjI
?����Y�A�@M��z��x���;gǒ����f蝎�+U�v�B�z9�n�E��cL`�;)�xWd`(�;�/yHw*n�]\��/�#f�J$i���0���Tb��b��!�3H?YBU[wt�'c�����Fx�%�
�H���E�ٵ{�����4���Jhl ����A��.��e��ĔAh�?���5
e�%�d� o�@T����6���v�E�.��Ap���dŜ�����Lm���B�+�;?H^��ރI�Hd������Г��u�k�Mvp{&;KE�A�ä́O�U�g����$��#�>D�1	�0��,~��PP���U�� 5wA�eg_��g�����߈U.�09�5`�J�p�".�!���*�d�/�$-�C�|�����O���û�P�TnQ�0A�tV�G��79��<�q��[�zg�qW�����o\�k��$(>_��U4��J�:�q(t�
��n�Do`����F�{���$�ri�����W?�9Q�Hb�"�m}�z�����CC�s��m'��(K$�\�]�q�oa� ����(G�b��K`�ۿ�)(�rֲ�Bm"� 5�P��E[+_3A�١!҉(	D`;�vہ�4���zРԮ��a��=����8���|cIb��|d�1~ӵ����Q\#�b����d:���UP��L���z{_ L#��TY�I�|̦�r�_D�b\w��g�3�$K�qf�2�K6x;9kT�-Ӏ]�ѡ���/a�O3�9��ك��]�Q�c�eK�p6�>�'�2�ܖ�E�o��R�[�d�&L�����F��,���@��⼚�c4�լ��Y~|7x'v@�UٳoA���n�������;�h���u��!���<��K�v�|�~�b8�S7��j���^k�Ŋ�s�Z)�@�zr*����U�l� �N3X�'��걹{ͺ�+�7��?N�ٖ������M���JԲ������U��gO�ԶB�p����#Y�'�5�0�kBK�n1ca�sԫ##/l��Bo��Ֆ8d�JL1`,�o�!�9Y�ֻ
�D�v*(�C�#�3׷yg�.��GߚNd��-W��JiVEK�d"�x
�M�V�ݘ �T;"� �pһ��6�屍��U�5��g��iϟ͜f��7:��@EQi���:���}�,m;6�KfG��b��@}�}~-&�?��Ϡ��Wҭ) 8��}�+ta%��@��JTݧ�{,Q�8Q��H�f�-�ӣ�Oޔ���T��Z}t�����`��1Bh���(�	6���(d��-�A�@�T�4��W�O4����a����0����"3i��Yl	%��G����W�l�CW�%�=����j�j��qwZ�IXP(��u��R)gqD���ed�!% 7���<݅��8ft������!J/lE&ư�O�3�2���OܿK$o�O�������bQ�_/g�5/�����C�_����Γ|�wq�46rZ+� lR��9�FE��m�l���B�����긕*�_���QlI� 1`�iSX��zƪl�j��MV
��:�~�PzR�[R��\B���9	<�=�
~�H��D���N�%0Ѿq,��l'Vz�"2wc�:�1�>̹)�^�`�L�p��+\���9��h�x��\���h���-�9*3+�́�U���P�YT~�b�íL�◛����b#z�ۊ��51K��+��R�u�R��kMV����Yb�Tl>_.�m��0�pX���/O�)�B�@!�δ �-���c���Hj�X�w�7A�W��������	{@'p"��F_-��Q�u���O;OŨ>&;�$��~�Co"��mC��G� O6�XQ3��u��!JAO1��
~J��~�ۺ��tn�4��
�)Er�e�!"��x�qj��T(���F����J*#v�4;�y?�ꏵ&�7�$�Xb���>E�(#��'��aB^�E�>�]
@����	�/]�R��� vd�sa����3��Kj�N�ձ�l��N;�����y���/�~��k���Mg,���8�_H��9�;����o�DC*�����:�۞z{����<�I�l�<��א���(��c�Vwr��\����3��a�[�Ɖ�E�g���j��Fr��K�F�l����u��oԊv�p���q�Ǫ�&X��`ȡ*���ᾖ��e�|Ou;C���w+�62"��BefM�r��cVBp���$��q��H�F_ފ�e��!�����E�IT�z`)쉁#���ؾ�k-H0)�_x�����s{}��-	N.f3l$N�iTD�d��Nz�aSk�V�w�=c�Ѿs@9�u���Ԋ�.@ �xS��y�7,t����^��"�O�Ȯ��LbN�m�����E��dV���6��Ǜ�-�9~����	�G�F�p���}������3՚������ �&e��R�H��h!����뉣��Ӕ��U'��r�ӊP]̯:��;�' h.���󷎲���)Y����Gc�û�\�"��s%-��!Ȼ!vZh/�F��,Dy-v��s ܼk֞�G���A���q[��\�wqn������WM���%�v�����Y6t����U�	}yG8Sx�(dK47J�i1�j����Ҹ��6�w��fC0f�a垦����=Ʌ�χ��Tx��\.w�ސښ��CWDQ�H�@�����1#i���\�tD'�m���ag&�Lៀw"��T�d�|s�T�7R���T�k}
��'C��jM�XA��x`�nnz�;Ա�te�ӗk?��}�f�cgpɂ\aw�9�1�v�-m��ͺ�������"1HN��7��!p�(�ҹ�2/D���Q���8� `QXH�@G�H��k���i�����G/3�w%�+�6��pF�h?������W�*0D�&x�'�s�:eH7=��ݣy�:Wt-�Ub���z���;f?����q�ٳڧ�5>A����쓽�<L��B�w���:_�f��v��,�И��c�e��m���S=_��]�Ү]��/E��,�)izs���6��hY�g$�#�ӯTc���JH̊���F�f����zb=��vym��
R�Z�Y������;�<�(�E�$�Wt*���."�Rx�C�rLf��lN�̝#Z�ػ=�M�҉-֭�fC�H���C��33�jtq�+�e-�Qgy|q�f�C�i7/۫sY��0|X���hw��Z@lh���~�o��{�綿K���!�~�Jp7�81^u�wJH-'���G�O�O�Z�!Q�Y��[�AT�E��Z[3:�%������L�bl��o]bO��J?)zw��*h�
��,	c0;��<}�"��ʪ�M�z�c�=��˺eW=�9~DWA�85SA�e���x�¤Q\�J�<�\tΉ^M�#$Gˁn"Vc��I~��#�52g��3#�������>�
&y̘f�P���|(r�s@����?���~W�*{&�]����B��d
@r�3��zX��?f!���\�߁z�+k{A> �:�7��SSH�>��u%�;X3�ʙ?��%���,ҥ�`y� J���Vb;t��1�q�:\��LJI���䳍�-Ipu��O���&��39"Gp�4N�DB���df3�k�r�M��K%��\��)XAU���\�R���wY�tp867�OGb�_�r㷈�1UG��P�<�q����Xo����M�_�(�~�Mq�yyd��؈�����8��U^�g����m����3��3� !)K�gT'�3E0��rm?��3
$�}i�yd��ĥ	���@�m�2,��>���n(��{9���[�����L<�E�K������1�y��&�G��"L�J0�wD`��{���4������(�"�h )��"����cd��i-��F�m�i����mG ܦ��#.��a�y�pE,cb4 x�� SA��7Ƈ? �<��)5�)�n�!x$��n{:��_�y8A<a�hl��!>�톍�ޙ.z0�o�	ŏ0������L�ǫNb����i��lDjۼ�ܐ�hK��	`��5a-�}�V8Щ�_��ǡ��xS t������$4О�,!ŝ���_�V]<($u��󽓅s"�I@����1`R}~�y��3�֯���i�9�H�?%��88y�1�noN]�5��[�ߛAH�A�=�UT�#KN�l�G �|E���QԡǨQu��e��c1�3ɵSBf<?&2�g0}+x	<l��VbĮ��ah�ꋆ��'��*"{A����u_*��dC����s(�[j�l����M���r�a�'@Dqs{ �N�܆��3�s�y _����UQ1�[�J	LD~��նӌ��O��i8�P"۵5S�U;~K�w��LW�����V_��B(�႑OzI�#�������:
q<��=;$�o����X�-��W;Y�4yrX#E�K8���������}�_e�`b��{��mk�Yͽ�!d������]9�O����N
�˓��E9��taR����S�ݢ=V}5
'{X�'�d{�m�=->ݜ�!?�q�0f FO�8��3Resd�;���h�F���
���;s����*&<�J�o�M�M?_5q��iN�����S�iH�b
�}6��??�f���֝`������%�f�`i
���٦�i�Z�%������?@l�z�%W7$.S�@a������l��ӆ�<�lZ��4��*������� 7H��UR��4�ݐ_E	s�@�3*UT4]��Vm�Hc�;�_Z?ҧ�!�yB����|Z�L�y������sN�\������b>�V��F	}E¦}��>�%�J^�_��{�Ζ���3�A�9�����T��R� s;*l��jܣ_���z�~��@X�ʡ�j��0ή(�S���׍�rDa�	'�0f�wSx4u���q,� ?(U�3���-�������n��B�c�3<���}t��E: �r+��}�GJ�>����H�-$�A�l#y��Y�Z���U�a)���^Y��'��"�'ID���mY�K2c���9d?'��&�.4 �Bipų�B��ke���[!Z>�&�>����>lD��#B��,ITdl��x:Qҟ�af��'��ji�õmr���Dr��p�%��%�=�~A��օ ���I��7i�Ӹ�[�Ҳ����K,ܽ�a4��[t��Fi.��j����M��s��k���Kl�'�J ��F�%L��"�Y%P� D|��m��N,��q`а{��$�|w�So�$��0�H{�o�t[��ҧ�Ժ	ǹ�o����4���-�Qgw�)2��CM���b>%q<�?o�s�r���v2�#_4�;�C�m�P�Y�b_`⺙�LV�>T��P'���v_����Vi��������"�H�E�g�����6\-��]�`��&\�#)�أ��뺟x�M�T&x!�/�	t>���y��IU�qd�3!�_uw^+�_[��V�oP��S��w�8�Ffӊ����zB�䬄��m��Mʻ.tw֊��0��SH����8�?�i�}��a�%�Ð%�'�g:��w,�r�������4*
��8���C����4���@x��`-I�c@�AYm>�៧��)<����u�*=�!7���� $�Ґ�K�m�pX�&%{Je�@�oɿ��%&�Z9�M
W����G����T���r�o�C���ҏ�+ޤr�E�A� ��u]�L�驡F��GD�zk��2�'Ш+ ��7SMfo�j�Z��JjޔD�X6A'�'��aċ���EQd�a�P�RX���\^t����k�[m�R�7���%��p��g�U��J�Z�	�N�[p���pg�m��_o�۾�L:}�Cb6���@	7�J��D�o;��09B]!�T�z9��S�~���E�3S����
k�vKR�=��p	{PF_��2�M%�чV�T����� �����Xd�H��i,��bP�x���6 �'s�V��>��Px�S�7�\қ�b3p^���eHo���1m���ǩ�+���m��_y�R�m�uN7k�n2��V����%k>����a^��Z��ZfѮ����R�e����kɐ�%�5�Tv ����)�d�n�/��^�f�O�b��(��Z@U��_9�x�����(����6|b�s
�;����r�U�)Y�(��i��O���,Z�9Ҡh#G�E"}�/@�7ys��*�5�^�_��D��s���,�2`b7�d��>O�Y�$�g�� j�
�������=�!��rr@T 0��09'y�)f3k�f]=�G�a�	Ȇ��*�*�/��ܻ�O$*�n�8�$"%�ZK���r�Lv�@�.���1RH��QT�H�n�jk&�%\j�;���̆���~n�9ק�X}���]�܁�Qtp����mW�G':���-W �8���1G\n��������B�j�/��jS�അ�j�gμK]``�E���e�;���mn!�n����߻�lI ���q�5G�0ޜgJH���8Z�@�Uj���:�p�ҥ7�����b9	cs�{F̓=!�_D{k�.�n҃��9�U��,{��~��[|��!*���:��a�
�9p��8�O3����0g��V=?y�J֔aC!M�:���T���˷����W������r(�bR�!�|����vf����Rf�+�?
����e�A�����MP�i��U��5��>lx��#��l���:�	��h��~���n@��̆�<vԌʮ�^��@�
�΅-k^K��E!6�{�iB}�$�p��>�\6�žp��f.Kǘ� _�����3��֣j�s-�.A��@���Јڝlg§K���s�Ղ�lA|���K{�-�|���4/_�(�RIevHYL��������w@�Y��h>]�o>��4:�9]^�͚FMUV����k�_j��]�)��cm> `������8���͹��VH{��
���N\E���/�o�v}G�k����$5g��q�~��I������	(\�
㊥���Y��"�y�t���?�ݵց��&�	��xW��%	����/2�I	�@J�ռ����Glo*Ӫ�N:ºǯ���[h�	����i�,� 5ڜ^�Su%�����KG5O7�@�M�q��%?�⠃�3��:�+�*5տ�݀�<)�����06,͇��y��)�	2�zD�͙tĲ��URn��z���Ҙ�P"��{*���n��|N�A�T�i2 ��&G{vq��y#�6�����ҧ�4W�KB���}I'������&�J��F�}�iP�
W�CF����A+�!9C�Թ�}�TN̷ֱ�n���[�Q�X��j��F	%,	=�ULJ��don�ɍ�ސ���E�K����?g��[#��`<���{���8�S�F_O/S�+@~�b�bm����(�ݲ_��,Fũ��P��qb�N#���n�t�h�"�p� D엄$��p0p���N�Ņ6��h9[aJ��k�~c>Kң1w3lie]���;��G%c��K�-NWM�Ӊcѓ!���o�&m��=N�߰���b�m���R3�n�D�G@Aj]bX1B�iŶ�e~NvȄ���S�?��O�/���޿S���(-v��w�H��M�$¢"QY��1L��˙T��Oz�,����;��y��ߑC�kU�SJ7�܁\4ae��E��"o�Y�'7�B:����D���Q(�jW��'N�z/��j�_։�p[]GPo�֡�D��A���j�J����De-�pTJ��*���	��o�����[��Ȓ�W���,jw�6 y!b��f/틕��vn�����[\��?��y>~�B��^#n�}�9�=:�o�ʖ'Hݫ����碄([EV���_s1�7�)z��Qz=�b��T��$b�����/Fv�(����Ĵ�1�(Jc���~�j�8��z�l%��G��
[G�5?�7���}�8j�/�e?�
�mJ��Kj�ҏۦJ���[3�&���r��!���3>�i#�$,�p��xm�^���Z����|�����s�����(���sQŚ��t=�A��<<���'�m�d�|[K�ḃ�ېvl����U��Gt,��@�)J>�p�>N��
����rr��t��O*h�-\�@{jNz1�-�=��밡���z����n=lb_M#%Vۑ�b�گ�)�מ J�0)m�S�k4FҊ���j�38�s�K�j�^����sX�u_�/�Ǣ܌�3�)�8�H�20+J�D/p��Jy.0hg��F����{��cQذ@q�:2�9gњR&��=�raD,�;�����>��&�C��Q��h�~\�l��QӞ*��7BFX4r�ţ��!�j_�L\C:?N鏹q�Vx�_�g�	
��Q�̿ڝW�' ��^E�����	)S"������Y0J$�lƬ��U=�\��݆<������`�Y�������4��B����H��Krń���;"A�H��.�����w ����*m?�ٛ�HW�gF�YF�})=�fw�2^��R�̖O`I�:�"���>L�.��G��Z����[
دa,D����Fe͡�,�3`��&�����gk�	h�N�y�`�B�5j���V�"ɍу��d ��S�n�I��&��ݫ_���S��B��Pv�~p�T F�%5���0axR�ۺBL���`��6Q�Th�y�2�bM�9�5�)�-',�),2,�}Tء�z�U��7ǉ�)*���rn�Z�jqE����Z�8(��+i�z�BUD{����ktTZ+�V�%G��Ò	�Z�f���ڒ�v�G�qآ���Q�u���[W@���~(�ӎŦ9���yԕ���D��lؽ�q�s8�K]aP���O$G4H/��p��F��<��i��rїM�fS@�4�cEho�(�ΜE�w���Un��ܶ���LЛj������w0�
�^]Q䱞��a���k0*��ͬ����"�r�n�s{=rc�b~��R�o�_� �l� �������O�@�z���=þ������~�櫟�9LM*0��;֣���vr4����m���k=�_W��;�o�t���v�McH�{S����8|"�^�(}.="7��8N�l�o�����psb[����c�"��v*�:W|a�Y(E����SЩă--���� "�	s�j�����3��1���r@v��%�I��fu�Ԥ+�����w�G�Q��D���	E"-�_@�IFy:"��C�B����Sz'%�_���<�7j����#-�K��o��z�Cc~~���H)�F֩r���}y���K�.��1��
��9���{�&D��q�0\��:q�P�Y�ҭmB���1Lb�]^�%��)��,����w�_�3̵d@��c���|�񥦘dp!k	��|�$f�ys��X��(��_���p\�=�Hh̆X�,`�>h����]e˱I6�s:��i�>Z�i�O�aH�ｖ}�2���q��d�Է�e�9@��HBF|3����c��ep�I�2>+\��^��j��� \%�Қ��,1�����$+���I�Õ$����]r��M��\J����70�
�$'�n#�lb�x<�)?�� `	Xk@d*��r�"�fI�A@��;�<pK�ֹ����Nѥ�p_�&z�pJ�$E�b�1}锖.|���Y�'!v�}�6:���l���_�qhe�=$��JwM������i���#h� 5RfjǈT���T:�G�T�(^V����l�UD�>h#�˪�~z�V( ]+�a���}�]���_�^K$�0ngL> T���@��[�t���c���L�Tn{�EU}�g���k�1^�Б�N��������~��ڟ>�R��R�j��X�*v��4r W%qk4��EV��u�R�R��L9�i	���ɱ�e�㛔�9W^�T�4�gD��������C s7VbK�B��%nZ�(*@'e�6i��%���?`? ��2�撯w�.l�p����L34U�]Z�Y�������N��F�3d�vob�F���ˠ2u����y���>6��SLa:����4%$�>�s���Z���0A0
Vm�?	��V( ��<f
n�Mj=�jV�nI��X���X�u���(qปد��� ӽ�@M)�9��Ȑ��ǐp�[t�?�uXA��܈�yk�X��z`��.�qR��aG>����%��F�|���09��J�/G=�.���~�5�_��v:���Q�&���ӷ��g�����1�'$v�P|�6�;����Tw����wy�wrABѐd�}���4��-��T���v;���H�#�Ja��7�@�}��L�E3A��1��c}�5{��Hܘ�hn�ݐY���Qz#]e�����$J��eڷs=���: c~%5��U���N����!�0�kn&���,�]�,b��.����N_��<�w��#D�`-�9�:r��3m�1�(;{Z�Z��9�JTa�K1��Rq8
��i"|ɻneͶM[����,oZ�����,7�#%���W���_^���o����l�U!�j��e�Frv�b��?�?�����zl�q��D�&��^��>��I��^Ye*;/�`}Y	4T�E
�"�hW-a��t�Τ���zN���>:��/�� T-.>2DS��w���/T����L�^�8�c&3���SAC�X�p����f�77psu� r0�,�8�6L�2��1а괓�_g&��K��8W�Q�'�4���h!��J��+@�Q�O�8L�3��I�et��,�wph2�\�#uM����ߤZRrlPr�ظ/z�2C�޶ț�׽0�R��9S[��Hΐy`��3��q�JGr�'W/v���Tv����ɇ�џF7Y</�Y� K��=�������Zu��EU�ڗ6m�[9��'V��~�9P����a)sа�����&���	̵b��C9���&�J�����Lڈt�YJu[���7�0w�m�˷z�$$�ˁT��8�? �}5��M}�~C�F�ֳ��P'q.�ʯ�P��a)3������~�L<�΄�T^?�3� VA1����W)��f��ʒ��3�1Y���d��.�#�ќ��,;0�5E��Q�Q�ĉ^�޴MO�~Y؇�%��E�1�3BR{��9�
C�d��8.�"��L�u�Y����֯�/�'������@�3����< �@ȋ�1���dAC�.�8�{��3}d	nԲ9�C�0h�KAm1�P1Π��#���"��~���Ba���u�⤠j{_�$�򱤴/��ـS�&}�@��EA��a 9{g54;�S0le�9g.I���"����eq��d�g�����'g�~�HK޲ךy��9�<�+��l��"��W/�Wڹ��1�S�fj>3-�h!��,~�.��k�LѢ�-΍���)��i�}�ޢg}/��Ms4~�K�,0����qM'wp�#��@�VQ�0�ӫ?p���L�� Aq�f�|��R\��@��/9@��E�ҀF���rB���Y���;�	�I=b�Suy�R�$T�W<QP� Aaq�]�1k�����._[�@���ѷ�*�L�!yg]����J����������a-�R�g�Û��{�n�8ս��u=c�)���m���w��`��!��õB}<+��Rϔ���{�q�3k��4�ö��Z�]#\	�4��`"���`��5��Z@�if7{\�rT��i����巂r�*�O3�����ks����A�L��7���4�O:����['2�)��:�,�h��!���=��6��p8Ǘ�W�ᖄ o�����R;l�*�O+yֶ�,夰\�O}-Lq���M��L�&w�� Yߖ��kÇ1���� $w�,��<�o�64��F�m�M�H�Y�@��of��Χ}�������Џ�~���*vՎ�,k��0��fwW���x�|�62�!Z�qJy��6� "��3��ڡx��O�h����'u���*+%K��ndQ
/�_;&1���މRÇ�/q�s��!�3#c��rՍKr������ѾA�9�Zi��;=���.$��g-�R�?��Qi11t�&��X� zyQ�b��$�<��*4�"�ma����f_y��X���@�8��Vk�؏qf.�Z?����0��-l*w�q�H���E�d�#��aL,�Jh�)�l�2�@$}|[-��M��Ď���C=��@�#Xs=��Ģz]��@9�}�\��+����9DT�J�Xr�ODw�K�?o�Z�=����L��l5`J�2�[xr���M&�.�/��J����(u �t�F*T �/�?����b�!�1�~�գ����lՃo��έ��'��4;2ξ��A�a��.�Ʃ[� D��K��ӆO_m-�	�<~ы�嫊��P�Ib��@lF9ude�m�����䚞#�o�b#8�d�%y4eA{A�vM�^//�d@�����R:�".��n������X���OJ^|搦�x��#{#Ϝ�#d�jӏD�a�
�6����0�L���lT*�l+����[�,���D�k�(W�A��N�;�W-k?`��H�&��ry2=+h A6�Wj����nga�O����b!g��O� ص�<�@B���$_�߶����rC�m��=�$�xA]~"�l0,Od򧅵��j�޾/~օ�Х'��n��E�|<r�7!������U�瀟��y�0����[a�)~�"�����x?6�&��zʸ����ä�B�����5�<ɢڲ�eb��;��Y�d�N�]�����U��F'�E�Gj/i@P����Qe��t��v�y,�p�&���-G^u���nPdX�iJ�X�v�y�^��E���5Ω�F�:�p�kHM<ߞ��Q��M���ųE:����Y�.1��)�4:�u}#��xCo�|�n1�Ҏ�{���6��7�=����t���L?5�U���7!0�)��fH�� ܻ��� y��1�	�DQ���gS϶��OEڅ� �4�i��1�-��ګK+؝x��g�P��X�/�;�������AM��{���륜� �Ĭ"u�R���,�wLPA��X�ɇ�r�h��D��~iPa�:�Bx��lGi:�u��;���x3BKz=�I��4t�#5j޵�����X��5��؋�	|0�m�T7��Y������CXTKU%�u�� ,Ȓ��Op:6%r��xf%b������]����#(kn�iJp"3�8i 8S��q*�4�@ 6U�8>����B��^�`rϗ]|�}��i�s����ê�@����]?�x;l��F�;�@��gpƸ��eʳ0Ѱ����e��wv-޹mm�.%@�5b��ZZ��,�� ��O����w*ǎ��=�%ѵ�c}#8��h��>T�쌊
d��&53?gj��}Z�u��^�|��3tq�#��FO���/�����^�(�%�f�d�k��¿b]�1
���W��#:�)�Sr�u�Kc�r�/�$.	(�(Y��]j@C_�q�ya�k��n��:��YvJ�q:A�	��
��/2������HvV�"��q�&���ʒT�JHAmߢ[}�Z�1��2�e[ѕ"C9M4X�yC��mNL<PE�&�CpCg�����۟](�A �<i��-���fJ��Y< `�zig�-y�[���t�p�B��e<�L����AɊIj;4�9��捉��k��d�=��<�����Q&m���{�^o�k2���e5O�vp��6�OL`���N�И�����c�{9�wK��N�H��_(3��Ve�=�`Nw�C����^�f6���׎w�G��6{�o
[kc��0�*��FSF���b[�e�p���ʘ뭈�I�lI|��C_k#��T8��e_k��ׅ����F�$�TF\$�o�Tbb�Q#wi�N�_G�=���cC������\,���CU����pZA��T�O[0ڕs�Af�:[
8�͂:��� ��A�E��a\�_�go������!���_֕��P�K[��Q�PGTj�Fh�Od���a2��^~to�X}�5]yK	�&�:o?�W"�E�u�]ͯ����~�F�¬����Lr�O�eQX<�Re;�/���� ��k�^<��wb5�]ȫ� ��,�z��q��	�s2y?k�� �QI�Ø�-��C�R?�
T^��@ǖm厨�%��a��EJ�i2)/x��T��T©�%�->Cϓ����c6U?MY�]^��H��&u\�~l#��Yp}t��՚5\���fs*�Bi�&�w~#���ō	b�`	{=�t��y���DQs�_r+�������WL�TZ�y6g���ʄB���+G+8���G��g`�A�_C��=�������b�h��[�$bJ,��3�\�3"/OC���b�[�Ӷ)�}���w�N�M�'�n�\�-�\X}o��Ic��hM>�(Ft�3Z�K՛,�0�k����{
�������/ۥ�۩N�v(2����kٛ��^�1��d��kJ�_�w+;%��Y�c���E�tGA�@P4B}n)gj <� H�f�@U]_s�,�R�����o���\�Fu��E?r�q'�;S���j��C]����X��ɝv uA��� �&�2 ��i� ��{ćB�֛j�Soh���Bw)�k�g~���-駚��	�4��O���afV�So�h�������B-U�GN���!5�cTgo42c�*�-8�;d|t)��h�6�8o�:	3�E_�����>���9���I����_�`��O�
:ԀƵ��vvI�=Tk�S<�ԁ3M*���Ӹv�h�&[^�3b�����N���%��=R�t2�t���]��Qި�gz���TG�����wu����9�4����?Ν�]n�������	 r_o[��x'�Qmq,��p�'���C��h�kk�$�H&����}}�nl�4_Щ�\�P�=�p%�4��	�����ĕ_�7�ڧ���A����G�B9<�8,Ӊ_�����qrb"g� 32�i���usLfN�����mC֟�Ve>��ْhB}h�K��Cqh�����ڪ�-,Yw���	�Q���s���f>b�Nޕ4zS���N�d�[m���T���A&.�ղeͻ�u�u�u��e�)�i}My`O�u��gr�����0734^�͢�:-�k�����bDh����A� ���V�(B������I�Fj ����ҏ�\A?�o&@��3h*l0T�� ���;R�<8��1�i��z�EZ���&�=?M��/�7
����� �3�SP��iĽz��]CNg��B��~�\������;���{MƧ�[���}�4��\@+���ڮ�=� �)γ�[�(�I�5/�q��c"�k�ڪ��2[nl]�!�4�~�Yƕ}MQ�g"�lrt�]	Y�Ӌ�Ħ$K��C9؃���������E����p���-�P/�l�w s��\��ͩD������ݗ�U�M���Uٺ\��?����SZ(?�/����z���<���L���%�o���o��^NUףP;P2��j�bGOP s^�%��Ӫ�	�tj̘�L�#V2���'�������|�/�.��0ғZ^\� �AL�{�`;��lN�X7$�� 0&C�R1�����-�=V.�r�t����G���+��c��#I�W<��l(:��?F|w��B@X�˝��������>;po�F�s|E/�0#(�cT_t�U I����}�0�^nN5jD��ٷn�w }��Gh#�Z�5esյ��Lj��N�Xu�?��U�̓�b�3����5׼�n58�[���O{��i6����MBE
�]eLm�� Fx��B��r	ح���C��^&��ĜG����	�vC[�y8Dg�_�ǿ:F>t�ɾ-~,�������u"���g���#�>���/���|��A�-�f�P��}K�$n_��Pٛ�μ����>�/��m���ȏ>ߌ���/������ڢ�w��j�V˩x�+4rs�o�.�O�! k��|���v0ktϑP��ô #m&�^�� �����/(����YRr-�{> <�-5q��&��w�}W�UH�n{�݉;�խ�Y�aO��X�KХl�Cl�����d|�u�U�G�)�E�
a���Lk�V�I����f�^�O�cDBB�c��X��;��cb�ہV��B�_��XoU3) X�N��U��-rz���ca��g�E���6��(�S��^���r��0�W��S�����h!�7�6�;�$�X{�b(���9&޹���$`	y&J_���4#��w��5UPs��jdJ)rR���M�`Ԋ����P���5��s"�WP�ig8�#+�|��OΧ.~���$�Dj�.��򭭫7Y�i��S�[��/ ���L{6�p|}R�����7�H&(6}OSo�*s��ů,����#� ��^|K�_�%��ii�[�gB��n�L`\F�.c[vޛ��]"t4G�]�2tK\�x�H\����Y�K�M�c���;w!�}��\�>��k"z�����m:E�(;��"N[w:杤-�X�����ԼE�����9��K8E򹰙<�,��S,%�vi���hqs�/缩�q�'h���(�|�Ӗ�6�`�N+Qm7�7|��%�ڃ˂���LnO�GHLz��TI�ZO����	h#�uwkЭJ�p�P�O��ӐG��m�V�`^��iXd�,�V�y�DW,�P���7�f�( �v��}�щͣ�2A�yk]qs�G�B����5�ڬ�����ŭ�v9�#5��W�,"vN�#�Ӫ}����;�h!僅$*Ɂ�}d������,����ѧSF��xk�X��Q:#��i;Csk����M�k�#d�M >�$\D��Ia6oϰ��S���S6�����D��0�2QЋl����Ba&�k�Y7JzoE��d��.a�zu���)r�/����E�_���j��J�=���pMa&������wՀ^\Pb(�m�7^%)h�|,]�a�wB���4Z��	�?X��"�,k��y����6���6Ґ�Я� ���X��o�����A��|�PyT(r�ָa��Sն�OE�/Y�+�Y��
ݏ �^gn7�+)���Pn������N�d��9GN������}�"3��*��j*���+vl8���I�kk��������=~`����j�~�]Sᬮ�~*�ꔠ��R��1 �^9�Z��7q�S�V3�'Ph%W�rT�t����34�LK��>-x�+�D�jf&|��cn��%TmE9כ�Uo�A�
��n�K +���,�!�Tsͥ�ʅ2�{2o��\�(w �3�CN�S���j��h�A�҄��I`��:,��yrm�b	b)g��@2E3D��_�K tg�̴���
h��8�z�aȹN
%#�[Zs(l�}N
��ݼj$	tc���$�z�zj�;4�a[���Zz�KR����J-kt�F4�h�Y`�9��bJ4�w�v��ך��M<��H`�F���o���y��D$�/�^Dl����͗��5J̫Y�8�xk��w��%3/D�Q�-'��n��P���IH9��P� �ܑ��J���{'?7!H��5�*����y����$��g��� q�z���~gr<̟����H�u�������v�DYn�0�u}#t��Qw�R����0OrP��"����F!%À��A���b����o�#ѢsC\S&�f�t<�٪qɩ�cc�!~m�/P�p�o���0�aw�6��kR�l�N� E]���S������FV�v�_��q��̜��]����;�� �Qz8�Pž���Q�L"���	����&�ֻ^�-����UkKa��Ɠq]�/�b��1�i��\H�]%�͜"�w�od?��eD���e,�yVhH.�~�J�h��ۦ�B�2����]�D�u�Z���X�i�.�9="�K�wm%�F����
�hUL��T
��D�R��P�+�l�#!Xm��;���Ce����� @��/�?`�FL�/Ժ��\`�8p�V�$:Ʈ��e��ə��r��d�N�C
�ʪ����5�F�3��&T\F_�Go3I�d��]񕒘��`p�L�-@��ln�dzrօWn�c)	���w��Zluu~�R7{����i�lH������ik~�z~o*�L���%�F�|������Q'cГ10e�.@��6�������L����W .�v�K?Gm���<�'�[., �}�����>7�=u��)01��/�# ՛6>�����2z�^mpB�{lqp��*t����މ�͡�w��>���������pBm��yn��s��T�}��]�>y�r�{�"��u`䛅/f�XLk^��e��>(u�6��e�����W
6�G������Ӽx�CVh��_R��9S	�p�u�,���*�?Ts�
�����Yw"Oo�i\����/Hh;ݹ7Q�'�TJI WWF"�PJ_�����|t��p��=\xF��\5	/�u!$�s�����n��J�(x��M�C(�[��G�L�����<����)���h��&�ٹ���)��$U���͸�\�?ˈ�!�&�2�㾲Mn>���J��#���' �A9�m�Z���\D}�JD���ƻc|��V����L��ţ�,������	�s��j�}���~J�������eO��B�=����_�	�b���rjC�5+�+�i�?����N��hz�wa��i�t3H}�ilϬx=�4y���ĝ�HG����Zb��S��e
[�w�?�K��՗�lD�1��'� ���J����
g���0V����L$�E�H���m x��j�ha$p��e��,�[m\�ZT��z�MG��?vt��{�	:�W* W��|[@�_�lj�]+=��0�J
%���*~�H%�g��-��KL�C}gvPڇdX��8��w �����q�W�i�(�-��8�3�H2�G�B�vAN�k��_�X��x���'���ߙ��du�2G�sZ��Yf�Z�|�6�,^]��8?�53����A!�i5�J�ctN2��6S� �"��r���i荺�uP����
�� }#��؈�����7�B����;��D_+U��z�H��)�k�}%+��?�B�p��Y����b=C��|�+���k1�V������ �m3٧ъ�\��_Żx,�xd��+�� �y���. �M����8I8�`�v��&�=F���v�
0�[<�s��yUee����	�q쳑�Hk��sC����9�U䡸�������� I[`��� �\IY^m����ږ�%a,Q�D�Z�W��r�u�f�X�.�V7����T0=��ˮ�v'+��LWNe;!��[���_�XB�Lކ eq��>��2n�͌Ps�����(�bq�n�}V~���?ƛrX���zݠ�,g�~�l'���{���O���)Ն	��*�W�t#�O�l�����R�NK�X|^lc����_׆�P��+7	=��Z���$:b3�F��Fb��J}�.�Pt��f¦�;cL6>�j�.E��:���$@�������BF���������{��P�?jי������[P�~�K���xa��U�S<�zg�T�m¦�ƌ'd�C@c^?̭����5���+M�?���ކ��q�K���ݹ�_CR�A�yw��e�ոQP�8x�~��r��
�T8��(���IRV�2��Y�]��<I4�LYӁ�pa�:}�2�C���3<t9�d�q1<�hS���w�	����苲n�3��t�#e~��v�Y^p{�R���-����z1�9	V������ɣ�������-��Km�MA �Q��WIc�]��H��8[�@�tN�р=5A^p����AΦ�N�ߍ�ht�-��yk��M<�P'Kb��p7���'�/m���s�[��W����6�`�'�ݧ��C�� b�s[�Z?�5?���K��\څP5ފށ̈�@/W�l���e��&D4�s@��c
4� �z~�/�>�p��g#��o�_t0�r��w���K�0*4��l6�6�_4d���+UΑ]�T�O+hA�*�����5��,���v��ho��Yg֣#Z��֪��ko�%4�/x糀�w��M�Jw.nɆ�����JA�`�]+� �8�.��jJ���^l�5j�߂6#̹�@�����q�"aG�������s��G���R���q�&>M�5<��a���������p��Ɏ#�Y]dSyr痭5��
ډ:Mp���s$�U�αكM��w�2s���=
���j���8{|[��&�ߎ�����1����Xn�wW�����m� +W��b��̧���E�L���@���8T��[/{�\�0C��|�I�q�A����qKҰ�o=���{�s�<%[�b���ՄB=�:n����^��U�d�Q*^mN/�r������T��N��h�f����e��vŨ�.�� �}��Ъ�zYe��R?`;����o���(� 	kQ�2��!�~��w�Ʊ�y8���|���	Fw��W_����-�`�R�&���-o���T#��<*��%�����:�u�-��m�oB"�fT�\��;xo
�Ղ,̅��Bԫ'���X�ۿ��`.k�5>8wX�$�����%�X�>23t��@I��w�t�O���GA˘Џ
�W^qKg^�f��=d��"K/Z�$|e�T�c�2���-�)��\Y�c�ʘ�kp�V!��/rtD~:p���*N�2�QI��oď�-A�^�	�V:�v!<�m��[}��v��W��G�$o���}������D#
s�lEMP�,��h��z���
�dK��xݬՋ��g#$)��g�W(C�����O�^�ӌ�/HVO��X�.�bZŵYT �櫠�P�����a>�� �{�V��<�*�Rz�Q|鿨T��^�'s���q
����Ā���NȕQbI:�V��N���������@qi�o��_ �Ѩ�mg�iY8�ZΓ(GH�m���?WR�~�qfui���	䄻Gkw��!�?�+���:�7}T���~���'l<��[��r ��zosL�un��~�T��*#��^8��s�6~�;J��J=�0G��j������^i5v�.Ҍ){�Κ��[]4��f�����	w!)3&�w���6!H�*�!�_�,B-�k$�c�\x����,���
�J·��7I�K��)�����asy�/��u_��>O�{NF7cPd�ڒ*vO���ȗ��ϩ	��
K�K�]����{����zͿ$xx��%΋Gc��df��wpǟ<���ه�^dc��� �k������hʁ������
��p,V�����Q83Hq��>Fdx��V
��q��`�Cgtv��}T���-��iC��"�ר�ra)���0�=k��rK�Y�����,6Y�L���|+1�ZJy�_��
?س^�aq����Y	�Y_�}yoZ�=��0�2z�(8T}�����>N��,��[�΍Y1��������1<ӗC`��ණV)n�\c>䮖wX���`S�,�����<�Zu�LE���{!�s!��)n�� �_��B���E�N
7b�d�լ%�CES�Ȱ�cQ5'�U��)�8X������Y�]��<��Hd,Ol+.Q��k�����E`ظ3���?z������� u�H��Ζ���h(?R��@���;i᫁_6�Y�f)�x�o�	��%�.W|ޥ�?�FI��F���+��Q�C�is)�.,`_=Q�x>'�9�s���yR�^�:����t�?��B�w�7Rt=��رcP��ֆ-<� ��-2�lF�e0��M��2��U�� q�|%PZ霔�1ƨ�S
!��V�'ub�d`��Ǩ'Zt�$k䁹�A�B��i������E��Ut�F�I�^-y��MF��)��S��RΗ����S^��9�[7䙬�I>E�O�FpE�X����	�xI_W�3��p�0�Y���Xc ��`#x q6ۡ�ٔ���P�O\����u՚JbOq5�4��z/U�Q���,�K��T�d&9jj\�w�E槫�&[�-�tg��n��;	�"(�1��q	��\�F"�a�]�Dd�)����ݖ\�nz���s
d��\�;=C�Ũ�ϝ�O*�m�"u���	����O�'O� �7`�y�Z�!,"<�Ѩ������N,�W�o�k���9\���k�� -��(��(G�����
�o�he��^�7�L{��Q�%���u��z9���pQ�D��9;T���UYn3+�&�d�UE�(G���`x�;M\Չ���
�D�M���3Dn�^�z��K*��E�ul'Z��2�����5I����o�fj��ȉ�B7(M��ML<`7Q�����/�J}t3�&�'IQB�4�|�ui9
S�/Ѣq���m9�ڂG
?��Tи���m��1���[pz�t��'�����+�.,]��!�@X�i���O�'<�z��$8}f�`�S���I
٩�Φ(�4'�s�I~*)2��lJ��"w�B~E/
���}��\|�F�������HVR��0׫��=���b�Y�3�Kt�*8]�\[OœC)B�t���_sVx�y�*����3j��a�nM�����흿{W���듰�f]^X| ��EN�6_��m!�C�p4�x7�B�B��,��F�!�a�n8P�Ku�JO���V��lڭI�K�L�oF�e�ixj�Н�5S�.�Wׅ��dVO0H��I���(��isX%Er^=R�Y���w��B���ۑ��ט�徬�<qIOיI �U���K�f�d �6I�Ҳy����47���uG�q|73�ƅ�D��SB�G�+lKj������m�x>`�������������/��x�` ���e�.������eǋ��"�T8ˠ�,���m|���;���p�<Ȱ5������S}�PT���0�6����{LJNM?3��9h�L\�����g�o��=.���d�x��l�wS�x�MCe,��H׵rUu�LH��ot�D��gy{d4��ʊ�����i���@<��i����#�
̰8��5��	��<&�u���48����4a;��ÿ����v����b���'gZd�Yt�Q���؞��>H9���V�9��<Z��@�i��(e�c�"0_�~��C^�JD嵺�K&�b���WA�@�Y�[�dCݗ��'~]d]pB�_b�@#i �и��f��+���XSŠ)����Z�r�a7)�	���_u�dK]�O<��U4Q��������=h�6�v��EX�
��5W^uFhI��(Gn WWL3\���<y/ө�  0���q����:�#iQ�ڽZ2Gb����L�|��Xf�zV!�d�� #�=-�Ay�p-b?3]>�����,������F��Hː���9^�ol���f�>^��+�Ļ�Rd����j,��,}�Se����%/)�����9������ʃ�A�����ڧ�ą>EX�` �P�)�ᨔ�;$�me��T�1e%�x:�M�˒�$S�z�c +Z�:@4d���®��	e�l���i���9a��߸�;?�yI��[�`����i�N7�>��; Q#�_	����.��$o�S�tk��Ͻ쭌���aoe,����^?S�h�/�ߛ�i�W|^#�;%B�����:0h.�,��R��!����FE�����(L��h��PV}����I]��#n����\W_?���߰ۜ,����]���|	m��3�ȶ+=��Ō=Z;��/B����)��Φ{h`NǸ�����q���h�XH��É.PJϣt�S�(;�^P۴��]__;�;`m
�W~���;��A��HA��dLP�܃�\,#��NV�J	ؗ��md7�V����0$6{�d���H�	ۃD��S8`;��
IvUF�@v�@oB�y�t�o]L18�ǃq�p�yv�nD�qy
7���t��!��RA���u.�ȍB�6�����&:\b���,�A��[��΍Pm!��r� ����e�HӘ�j8�����J4���@���O�e�9�����R�����L�	�Zq5�cǧ�n����D��� I2gc���Q��;r�鱹px���pM�ln�t���Ie�?�6���~'qW�i	$�.-��5�σ�q*+�W;{BD0��x�X���lNa>H"x&��"{� ~Ҝv�^k��Eӌq��%'��s��m����r�a^�beZ&��4��(+�ʽ����L��̑�د�/�/B���P�\��%K��w��bl���JFy����iBht7��qc�)�x]��ԷC�T3��S�`���$��œlf�F��� �;��r~-�D���g}�t�L�zgvEĖe ���ü��g	�%��\5ݛ�%5�j�D��	��㟷���]P�U�T�#�g6q��q��!������ͭ��Ǣ6�_֛�+�.���9)���2���F� d����YTT�3�}B�6j��*��\~Z$_��p|�B:B���5�����[�+ߴ�� �\��=m�?�T/T�a���˺����a���zv���18��s�rL�(]���|g������ح)�l}0֒Ǘ>�;��(մ��0r]�6|�̌�½��UIK3 ;h�X� r*�I�<\v
��h�a���
!��qI��t=�و,r?rA����G�/G� �È�L�s���������<p�!�U�s�.���jce5vi�e~�A��d�K��t��u#�S�&jw��_
S�co��I��r�Qu���s���;�����rMC7W�2X��v�tC��d�4��zqcĊV��x���?��5ɢ>*m��LUby	�	�)��������P�mz���l않ؘ�7��A��@�^"��IYW��3���>����f�P@�Tǡ"f�
���r͟e�����!���?����h9�(@��D62�A��i�_��a"ׁUhcM�)�s+<�/�u��S%����ɱ�8��;cY��m�б?h��ͤ�������T�Y,B0`�0>�@����~K�[:,��yɮn�]�*ho��7���32�$��`�#�*i��N6�#�f��#�8��&�t-v�:��bA���F8�75\�?��J��V��-����۠\�<���>�E�56_�Q<���Äc��ݝ����[\}��
�9[���yg��.^�,��e 9���v��X��F�ξ�~q���N)}�f��)u�|s�S.�ܙ/<_�lmd�*A��݅̈́o������[���A*�����W�M;�}�%Y�
xi�CH2��j4B2w��6{��KX�h)�����k�z���bsd���W��o�CYP����b�L�:���1�h���^���3�f�#V���F�Y��=}�^,6V4n�����PX�ެ�{�d�]�K��b�
�e� ���A�>Id{-,�&��������eǽ�,�_NʅTp����~�_��-ASY��.A��=��X�>��ʏM�O<�X�@�2VB������2��L���V�C3"-<V�T�IgBs��6d%�,H��6��A��@b�'d��J#۳��j4Mdot9�sL����mQQ6J�Xs�U/8��;bz�i��Y�ݖ�ݙ8�U1I��d�$"��ρ����f�C�b���D���B�J@��2��έ�9 tD�0CسI����l�b/M󣥇=���:�MZt6's%���¼�~�o��w��~3�͇j���QЈ�������=���ug�6~7��M~�?%���)e'��hq��MzNQ���K�Х��;_D��u�����I����7!r��فw֯�2QE�!\�ӗ����UMbG2���.���|#������ �>l�o��[�?�)��l��_`����V���rv/�nG֮��d:R+����};���l�v��z�s�[�ͽ��	�����ϳYd��Q�/j:L���6.	$�%]P�g�z�̽_3g"z<��?�Z�_����|�����g�?r7隔v��G^3���mo"n,\���HQ_)b'Φ����2-�����5��t΄d$�<���b��Ⴭ��,[>'	��N���Z�5Vd1�=��s��0-�'����<|}5�-�'i���b��y��/T"	'�0�6�Mպ��r�jv��r;�@��eR������wK���Jh��G�ܹ��>�V��1�'H���)V�8�$��������F���x�I����ZL���m=���#в��� 锾V1V���
��ɇ�9+T�h����k4��7�o�l�Fu��s�:;�&zA��ރ^���3(��qЇ�"]��0�{��ޅ�4� gh��F��f���1�Y�Ly��l{����6���C*��b��7XQfy����!��5���Y�37�~~��.�tj:��1���>�:1]7R�X�jE��c	�Ky�\����^�8�GRFI��RE��T7��A�g�N�.߽$�[�`��|B�Q�T�[%ٵ���h&n�����J�
d�!e�3;�t8�y�ku���,C["v�;){K~�.��>�8FLӅ��.M
�����Au�%f}$�/��/y�����A>���7���t�VT��"��6I��`}O�T���Ǳ��V������+�I�ly;E#G(i]U�/`�͌��C���������v���~`�7Z3vD��T�*�g����Ί�;�WQ���S������p}|�O����9ƞ���[c���#U�I���ć�`���N�G�Ծ���,+���+A�G
��O;��� a��.]"Qb�㒝إ���3����;�����!��N��e���#�K����k.`X�������oȷ�t�*�����c��|�]{�f}B��͹���[wlI 1�����d�e�܀�-�FS�H�i"2����r0Ǥ��~�J�r�C�)��h�H�g�._����nR��e����$x)*�q9��N~@* ��GgsQa7�`)�$���$C�./��+~�]��Ʊ��xC�W�VCY�.�����c3W������'v�� �+�5	��#,mӻ=�����:�p��9�� ��\QzF��E^5VB�b/T��J���<P�<1�e`�V&�D�[T�5�1�Z��*j����с��z���K����:����hD:�E�>>��1��~�O����V���/�J5��#�|�WU�a����fq����D�3��/�8k�P��Aʌ<%L�.�-��x֌l�b�����O��q)o�����*�G���G&5+T��Ё;�Z���0t)�tx�!��t/�Qm9c:�x�����̬�X�ؽ^�\�A�ۛ��JE1rz�ʅ��g�����۵��3��3���%��u����'먮�j%MD<&JEd�lyt�.�	O���{��΂�=�3 w^�S=��sR�J4��M�	��dصL�h���{͐7c޷jLX�?.�V܉s�wR�x�u�5�f�%�d�U��q��X[�Ǔ/"��{p'bH�cV=C���G�t�#+k��E�/ ��I��}(�m�.�d
 �v,2�p��>�bT	�;��#�5Ȋ�Azl%�s�`�\�|�w��8.k���G�mV�7Q�
�A�|���(��6<C$�4apɶ�A�o6"p�E������wK�-Wp���5y��=۵"��E@�l�h#�A�l��T�{� 붶ZL4�q?(�����9�d�_�I����Y9�§��y�g3Ѿ8R܉r;!V���{��)��`�*dd�7���էC]���D��Àp��3{
ٶ��JX?x�
\�^f\���' ]I��]�錊{��:��g��yִ]��� }�k[��R�q�(@:��4�q����q�db;���Y+,��h1A�o���4�O�����E�`�����\��&�{��aq%Z��������� �Z8,������ٍ(���E F8�x��gh��gFvv<!Ͷ�'*VY�W&V�[��z��RH���ݽ�v5��éh�{\�%���UY������9S�weH����S��>93yU��]�j���u��,34Ҟ����W��&�"�J_9��X/,=lG��Z�	b�8f��EX���"!K�����lʫ6m��<�11���I[I�;q헣|�����������p��w3�iX�Ov`Z	�m�V��|����h��AT�(�9T���a�wسw|�{��S��|'��#̃!�`�!@��Y�O�y5��5��!-yw�t�c�(,��A9�$�'΋�C8?��(s�sZa��,�1WT��T(������νFg��&6�
=g�U�
�:i��T���ۼQSj)��6E�.�G�g	"��Qv��4�Uak��ְ�GΖ��������T��
�x*am�ߩ�A���T��U�r��%I�1/tn��ڐ�"U`�a��3�l7�4�HC���[x.8SJ��O�s��Z��t@�5	�|8	�� ���N˒��.�K�!D峌�"@�+@���;�ʓ�|�_W>&1���t����q�ͱ'5�9BpY���_L�k˄?;�Z�y�6�n����
�ݰ� ��e��W1�K�@x	/���<8��Pdk���%_H˺O?��J6*�P��3XQ�	cм�<fӗ�c���h�4���Z#yC ��z��qbR��P'�?I��>ˇ������@�]����ǛSt�B����{����ʧ��uAy�ԕ�хJ��\v0���4�>5��B�4y8YA�ܛ� �dza�C�h���ԇ��4��OC��pٖVT��_����*	Sn������%:N��Ԙ�T�j�E L�2Y
h����.Ԭ<n �b<%$�5����߹g�X�
�4LJ��=����4�^����Mʂ�I��W��B ���{AG쏋
�b[��Ψ/�@{A]Կ%If��ە��y�W�J8h���fd�")x̚A�ҫW��.�����!��i2���u�����P� �0^�N�Q���iP+�+(��] �K�~EZ��ŗ���Xy�[$Ɯ�;Ko� ��~EL�ge��]w��e����"���+�1y�?�JDn�Z��W��xײ�.�B@A���u�ʜ$Eo,R��f!~]O�Ë��60�^�6g
�Z��H;(^������� 88W��P'�F�!õ ��cչ���e��mrt�M��n��t�.&����BY�@�.a�,�-3�[�qv�r�������t�a�Jy�+G�_
����Z#��"�H�̈Ҥa��䬐�s�4�v���R�#�C�:	�^|擸̘�yjm,;$)m���V�x��X�Kt:Ke U��˰�ж��*VD�h'4	�7G����P������_:��"\�eN���HD!�
���y���\G���1�J�m��!\�9c��w(QU���A<��e"���Cya��5�ߋ�O���%�
��.��o���ӡ���⠼���m�a� �7�Z�A�-���#7r��]�z\vRH�Wg��Q��ʄOckG�F��EO�ٳ�Ph�r���kj���#2}�:�/�����pwb�~�)@ӣ��}ü~ТEo����T���bx`��G%+���s���-�7Z+�C��-����7��F�<����
�tˠf�JݖT�wOL�F��ʇ��r��n���w��:|�@[�K���{�Z��ݡ���jEO��|U�C%����gx/-x{�@�0q�e6�,����QD�@}^!U�l�����D��	c_p��F?m�9���пX�͜�K7���)�l��αϵ�PS	�co���id`���{�e��"A�9! �;��$6�3�����W��^M��R�Ź ��*萮�o�S�A$8�o��������:�I��z�������s�V�;��tm��?/b*��)�+�����9�O��*�W����V���K�#�HF�%wk&�m�x��D�OH��i��� ��]q�)S���d�׭�CL�����G+X�S�#��;��Jj�`���f�3z�� )]�a��H������h�k�x��LX��ݱ(�&�M'/R�
/½�HtR���-�A��?�z�,���>�lB$e��K��lJJ��MMdL㛶���З�cz��h8{�N�r+�99�)�0���J� Y���=PuS;S�V�A����[A����ޟ�K ��t0��+pb�0��eW*�B�R���9�h�E�lŜ���K^�=��=	6�o��9Ί�C����簡�_��ܠ�t��Rgy8h�58�����FXƺ1�����\��~V�zb��}����Z��{�9���������AM�>�D���)C�J�i�	�U<����֙A�yY C�)��o�C�fn.^�NDG���o���͖�t9V�BD�I��*��1}i�pѮENnZ'�}y�CK⬠7�QA��d�f+�^L���$�h�ϲ����	�8�퍑[/���qR/����А����#��L���v�pgl|%9�g��Ky�~��O%�)�T\,���OL���8��z����$��E?��	I`��涘x�x�ql�;I���FE�p_�L����[cWhe�4p���/Ρ4U GД�ㆄ�����q����R8�+M�����;xI�Oy��-�C�/Ņ�*�A����t����Ho}���]�\((ta�2R�����9��.�����= ��P��I��s�?`�i���Q^�߆V��1��Ɉ҉D��m�tb���K��M���=	ē�O�iAX��O8̩�r�(�_����(��ǹ���&M?*Ob��.�W�xJ:Ȁ��HQn|��Y�d�Ug��H�#�jF�1��ޮ����!`���i�5���� �Sc`��q=�#���t)>��j�Ȕ�_��E��뢣�� !��P�ORP�d�P��W��Yj��2��Q��?B^Ñ�3
w�a�Q�D D4�Z����v䭐Vl�_�y�)�i�W0Z��nRg�3b3_���c.��[��h���k	�Ȃsm�o����q�ub��)������F5��B����)�h�ňa}>�w��)+�NYZh�7�JmM��W�\���~�Wؼ���D��BRa�W#č�)��z%A������E��=���6{)���J�]BF�W�[
m'���f'K)��$-U�e�0M���-|q�����7H'�td��������*n�aK�9�1���G^�ٶ�� ;~���y*>
�^+p8�Ks���f$�*;���o�v���I�rDb;�¡Q6��s4��.�������9rF�o�#�V�������͈� :�`����BFM@/	c�q�8X�~+<~Z�Qo�� �\32r� 6�ɟ��Bz��w�2;r���7��p��q>�T#W�ۤ�m"���	�.Ï~����������_������&��I����������cH�M�]�#S��0M��b�8�Y��2����+mj6�TϹ��ԣ�p�,�3
��	������P~�%��J�a�|��f�j���$N��n�뮟ɋ�KY��A%)IZ�����!�������/q��.����۪�٣�U�}���3b����q���dǒ����q��5Cj��M/�4$y��-�!砨�}�V�N}�B��Sږ�����6,�ra	�H����#c`��.��H�cj�o�F�'����~<1���jD������,��\!p�-����,z>dy��21��_Js���a�p�����m3Q��>t=1��1�eƳ��V�1�QyH�F��:�S�Y���󵲽@켯%sa)�����M�}"X]�L����孙��`�Z�V./PoЃ8����V����W8Bڠ�Ϻ0y��<0x�#_�����m���F� �5"aE��m]'��bp-����J*.-�u�M>�����C�p_(@���V�V�����⽨�ɶrЇ�(1�(!�iUc�{ӵ�-���n�$�h;�i59���;LQ�����Yߦ/��W���r6 ����z%t�����n�5D^����%�T�D��#Ҳ���e�:�;�&�>T����E���b���X�������R~QГ˪X*&�R�Wfur4���u�ԍAGK_����u(�oG5lT��ōI�����M�^�x�l2;�T��J̆�>��_ԃ�"��[BӲ�{Ѓ.�_F�8�Q��R��K�0�3�5a�����+�m!�iV�����t�F�?QI�M!���ܪ����뺦���O)~��^�Ԩd*뿀���CI7\X��O0z���ɴ[���%7E��\4:�7�&��<@O�}W�j
��Ę�¦ju)�n�(����26$f8�ֶ>М�mm�V�^o:�ڒ��W�e�����[њبի��8�f��񸟇_�;�� �:k��S��J��y.�ɋǥ݅_x2��*n�k	������^�����y̯� ܇��*j�lV��G�d�	J�y�S��v��W=V?aƈ� �%�n\�F���^^8��X>�n�:F�V��$�U�1�L�b�a��fP����f3�~�J��w�7�#���a�ȃ��R�ӄ�c��ۚC�e39����o�s0KAKA�H�PS����ӕ�ٞ��E�C�J�¬��E��k��Y�xx���vH$�.l�t��rZ�d�5��:!�S\�b��$ �!�_H�o++�z��d7��d��~	g�F�?E�?�Ԭ��� Ҷ�3��i���m)����K�4Y���T�!��@��<0޿K���謦N0Řw>&{S/w3]�-�0άI-H;w&k�%���}���Q�Q�
&�%I)�*du���})U��}�u�D�82���c/�w7ï[�㯘�O��(���S���&Z�C���+�3�?t��M���6�D�1�|m$q�X�I�E"��-H�����hE�^�XB"�,�_��og0[_�HW��ġ:�T��~�V���#�yw�#á���/��g�z�����~/Sjǈ[����_�;İrH�Y�A(�թ/�Z��&.{���xv�oC�N!-�J�84y���@Y{+f���[o����a�ϠQ��2�4��ַ��O	�N�*���V>�*�hVu�e����`�\�p�����y�����x�=�>���Ί�&��ޔ�|%�>�X��#y:1)�j΂+=I��/	.�p�DؼYݥ[���86c�|����0v)��� ��,R}(�S]ֺ�qp�՚���Z�dt%y��8�7��s�E6��)�y�^P�m���i��yyӬަk��m.vKE륫-���sL�1Ǘ�&,��( pd�"���v�y���3+��	:�|䐑�u��ݩ�Po�e{R��ϯo
����t�k�/�h��fRE372�2�ˉ�0�wx�gn!"/sJʲ��(��.��d�
փ4ҳ@/�ttŦc�~V�?����C�ٜ�/��`���lY���A�v��VYC/��L"W���%��/_��6���_��t|��mR`���- I��9K�}���[���Ģa�Ů|�����";�GO�Ć�^@~~��*�e��9�C�� 瞅sh_M�P��N��oLL����*����p2\A.H���j�QPר|b[0W04���kƢ������Їg�� ������˞�u��!���Y\�9@�q�qr�׸ITZH/}�#�ZD7y�E"jJ�Hְ���W+�3��ǹ�~sg��V*3����ߦV@d���uy���G���q�D1��������
%��n-���Y�?E���WM�)s�4��N��0-�ea�*�4��DY`[����\ �w�pӤ��&�ֱ��Z�C&�@o<bVc���k`�`�;��.�:V�p��<���]�pϑ�^z��MH�w؟}S��sjIU��R7$�j uz����\�0i��/}K�r*X1�c��%�Ơ  d�'}�|�:��`_��	Nx$#s���3U�V,�d>v��w%���>���(��&Ea��@B���]@�.�������,p�a����%��
��@��D����)CaN�*L\͓ѣ[����
���}uEfK?se�+LXT�#׍6.%�VE�>�:0A�Wd�����c��j��\������C��n)$%#�jȄ�-�!��?�O�'��rt.vl����ٛ�лr�~3��&r�+�q��ViB-��N)��T?��=�*��~H���������!<^�Y��~�n�6%�	8�P��ƙ��XE�!���C�"5�GY%�EoN��T��H�!.r�e=����r��uQ��j*MQ��wO�_�_����o��O�o�k5[3�җ���.�\r�O �`�Y��?�;~6c0ס�j�܏�vx�tQdz�E,F�ЎΎ�p���-����;,H<dR(�1K���i�7G�z�k�V����G^�w��w�hQb���A���C������y���P���E�6�ժ5�Q�e��
�.(~|s�B�����Pʝ^gIU$;�� �ם���C ���ouh�iTֳ�K��ARܜl��κ~������J-�s���,�'qM��e����n�,���wC!D3J���a�щ�$fW��A;�P��+m�Ah|���l�N��E|Ć�y{Qs�`��)ޞȚF�x�p ���w�����T����F|Jf`M���ʅsh�����3.Ah�����������V����k�?
�o��P�H|�>@���^�v��?Y-���]��x K����X���v'�뢓ii&�<~Z[\��'��lx5�/K�����c�XQ�-'n5C��,��a�%����u3�,�M+)w��Õq���nyO,�žw/��5���/x�� ���@ݮ�Ba8�pǿ�}j9��9?�B��?�q\?��y���~Ýg�N���=�=�Y��ݑ~O���t���+(�1 {�#`�������,n��� g�?Q"�aF���kT4-t3� j\�������ĩ�'XI���F�Sdǯ�e�5�7HK���.�B����y�>�zD3����sjZzߤ����%.q�I���1T��֤D	]�Dj������J�����#�Έ��2FYc� 7vq�:v�]ѿ��jy��/��{��F�5Y��&ot���
R�X����H�Ĵi[�(��|p��[�h%1�yh'��a�y�������}�C�G�b���68�B�d�̣p�xF1z{�T��*C�����h�K����6^_�4TI|:�5�(���̧�f��zB�ݏC@-y�Xy�?�q�N^�"~�ػ�{p����*��Kk\�@���dT�����"�תSX}+�3�|�1#?c��qh������]��A(A�+�ry �����&M|�`#��r���'�����)V��Ꝼ���#wݨ�KPn���'a�I��X/�䧓�!X�-�"g�O��\@�,�7E���y�-�A@/�c}/~n���J�O"9O�����U1�A/�/�ݧ��®�i��b�t�fV�M�FjS��s�lW�sZ�E���QA�#��c�e&Z6�y;��Fw��m=_�z���4�����1��\ �Nl��m�;M�A��)����[P𯵒��,��sN���-S0I{�U$�ԤLїl��^��(��'Ȝ�)'wQ6Vz�sZ֣YCY��(�I��KT�y4.�r���Ƹ,�Q��)3�a�3|�����@2���B�8��]�AXjO�4 �b�>���9!�b��f���g穏H - cړ��1dj?��:i����СJɪ�����o)d����Dg��~|���_k��}�?�gt�$5�eQx����&2]a�'|�ٷth\1�ʆ}�Fۖ��u�[��'�(I�P���x[�f�fIuڟUN�����]�eӏ�맛���a	2*\`�����#�~9�9j�hwp?b�D,^���}b��$=�Q!� ��h�<tbFX��/��%cy��p ���$TjH�IVVH�P���t;�ÛqGVZ<Ǥ�;����b�#�Mi��z.��+Ԥ�|�	�84���l�lT����x���pB0�m3Mv���=�QyXd��q)P�'L�8��H`��`W0F���!S�s
�>.�"/Ȍ$��N~�b@����/���ֹ�{}A7Clϣ!a[�I��ZCJZ6����x}��=i���鶩�P���ݒ������=p~�C�o���Hb�v�F|Xi$����Yk�1�.{R?k��at� x���ys**ǹ�ƕ�W�kq�|�G����g/ܑ�:t���}�+b+j]�>��0�h��g�p11�,��4�J)�ϵ�M�dn�~�������KR4�����-�J�XK�w ��shғ������A�ޔ����M4�BxT��;v~�)RYʌ�B���⤬f��'D3כ}��U1N�\+��ETZ��� ��ϖS�V��6����l������_��9�N�'	�v�H�B�>�F���D�gDZ��
{u��O���%��E��.�{�	�������I�>��<������((6틹s/�2՛�6¬��H���É�����{O�+t�*�m��6ȸ���;��FQ��<at��� ��J�I��_Á�WSCV���7�2Z{i��:Ź��;��b��]���n�7�^ (J*y�XO�YPq�X޳��2u��Ą���
KTE��^$Pw���.�d�q�6�/-�o+�C�(tU�m�	S�n�^ڗDG�6��]�"���t�{������}P�ד�?հ+�oT��x�e��f,�t�a��o���h@=T�;�$��?dzk��)�j�����m7S��5;������	�޿�t�蝑���L7J��}���Gc/2�Մ��{����/!��O����y�lXNB�xtb���5�jl3���,u�ȼ��FGg������8��޲ij���������M&�6����U �@�͚Bs���I������Yֽ%%����ҙT4'�X�k�ivrE��Q�7^�?D�l�K���_�Y��n��x�(����K㵱���Ӕ���KA�L*�x5��pL4���F�&g���݊6ȟg Y>��ճ��n�Y���-�5IK�)X�2M���=	�|BU�!�}'��g�1��׿6�u>c��)�4�B�$<'/b��u�ʃ�K�r,oF�g��8~��m�0"W>�,��͎]f�n�+�(�2�@8��i[=���WPK^��W#Mp�p�j-��Qm���z�EH��g�A�a���*�PL�X^�֯%LY����x�� ؽ����r֘�_�U@�п�dD2;&�q}�i�Q�*?ZAu�!<�����0=�����a
���N4x�v�/~��!.$4�>In/Ѩ��8�D@T��#�C#S=.�y�@�U��g��m�VK���F9Oɢ8-�A�Ğ6M`uQ̂K��_����b����=�$�y��K���&,]2��>���'�_G�g+Yms���A�:���t��^�_���U;\��ND�����:�cL���e���f��2	�JJ��lga��]dcmׅ!��5��^v.�!d�Ӊ�ފ�����Ĩ�[ܬ
S�
�9�|<�\:��#�����BB�A�p2+�G*�<W��^E�w���b[5񻴺�����-�DЯ�T@�f��ra|�� +��� �H����$Cn{S٣�w`��E*a�f?�^��b�W�j��G�A]EI�qe����8i(	ķLso�Ln�{Qn�C˧:@A@�'ʳMF�z �`o���ҥU�,~�M����2�]��W풽�#k��| `VH\���bS�ܪ�B��%�D+���-����.�!{��	t��(��h��ZX�1[�z�b>�a��nRSR���1cB�f&�=�]Z+�&�)��<��O��Յ��\B�I��/ih��1�%�_%��hX��n�V���T�n"S�2��fQ�[�8����A�Ġ��>�<H�.-��/O�C,I�����\�'ў�NQ�{4��P7h:�LR�aԚ �%�FҔ��tՈ�)���`���w�1�Y�����wGo8#|�Yz�>6,[٧N�s"� EkVo�CNe�9D9����GN��9]r䑽4����S�S8y����[/'����GT�+�"�����1	A�����/>t�G�1p�U�"���X'��AA!��9H4n����U?�o~v��*J�RY7+��re=qo�U�_���a�"T'EbГ���*3���b+� ܯ�K8(Ȝ� �|e�����˔㠇�c��'��N��
! " ���qK���[鐼�<dy֬i���)����D�p���s��������L��������:������]m���K&�W����B���3&*���z�K�y:���`���CGa5ؔ�䠿���Ŝ�]g���a��6���T,!8���@<EF� �;�	���\ÕoK�èR�А �_$�b�K�y�!>�
��UjDu�����z��&W�JG����:��}Uqfc�7���.����fH3���8�B���hu�[���2�j�Ь�3�NA���2f��UR��1�;py��؟q�T~��نQxp�ű<��A��՚�A�vB"rN��6b@�Q�[*��%��p�r$dHk��{�<*;���O��
a��>��>��x�Z^��"������7����`�P<����&&0C1e�µ��i��hG���l�}��ո['�1�^D�W!�ITl��X��n�d͒˳�%�t�/c��LF��{�t��y��yU�T��a��x��'ZX�U>V��!�x�a�tRc�����[��1���Zar�K�"���j�Mkkи� ;!h�mSo���{��Ęȿ��ԇA�r��"����:�2.%��g0K��v�0i}����-�X�?����X#�΁��7��=¸ޢ��y�3�|0��k����nw�zŁ�.eK��A�R�}�6�y������9/_��qnut�!�x|�����=CI9�:��Ӵ���;�|�g��3��:A���O��4���q��+�.�|p�K����Wد�L�l�!Z3C=v�C!�L�=�*���sP����d.�xc6AΤݹ�rLV�1��,�����1N��³�L�}�z_���_y䝧ǫ���t�S~���xYլ�Y�	F�����f vn��8�~M?�j�-����D3�Ac�p��b~K��rje+�|�m�J� Ҁ� �8F <�4[�'�,\�([ �Ę8���&6X��+���1*��"��!���CA�M������`��-FV�NG�h��_�}��ň燪�/y�HHQY&4rG�b�J-�Cz��m�)�m�x�yk.k"���lU��^f���=����a����H��C�]��i�$���`�ʌm�XL{�Ʀ�n��~ۅ�̣~r}?��b��X��?�	�d�'���r�7�X(Dn�m�4~��6&ŀZ�s��+�S��a�(�gC��}6v�kƗ8ɢ��M�
����ఇs1F�o_Q����9�����"��� �-��G�Җ�����F��Y��
:V#$�����C#�bLۀ����񯯧0>و��K�Xd�Lw���'A����#�Uqu�m��-#ם�w�;�O�r"��U^�";��Wh]���7�RN)��q`=����g���^&!V!V��dKp�zV�g!P
�M݀��.zq�Ϲ5j#�L	J�S���FoK�6}��C�[fwN8(I��ūH�"h��H�,X���]���e�/$��J	2�D�[��[r�E�q��T���6^O�x�!��ͽE_�c��7a�U��WѸ��FL���f>#��p%r��������9���WL�you~����D��c��p��e�9���Ѓ�@xk�[�g��%!Ї#ŝg�UHa�aR��)����=Ԥmt��2��S���6˩�R_ڲ��:?_��ECE��7��,�]�E�]��`�oZ��IK"��Q�`��<��D�l��������]�*������D�v_�JoHZT�[S^�@1�Fd�����&�f�������K6��~S�X!��{G�yON��Pȭs����<������m�JNV�P�"� >�	3��.*?���� Z(��dI�d��g8��zn�t�j}XlO���l�PQ~*8�ճ?��Q.��y�u���0�`:�Q
�e���@NX�1kPk��Y�!9��9�K�U�ʱ&!������I(���ә���A�.��7a�dqj��9q��Z�O�@ $�$'Ѕ��Aj�h��p4Ⱦ�̎�Q��Qg�.�48ď{��k�e����L<�8}�)/]���O�ㅨ���b�=S�qsT��"�J[����L��fRߡ%�� �]��>`wSW}��s��G��P
����!�e�/����&Lو&[l�[�y�s��«���g�r�Di����__Y��٥(�LD�Fm�c��l�Yf$Sq���u؁������7��.��-��WS��sx���[�z��Nk��)N8�|�Td�+�j�I��*I�$*�C�[�5-�

�k��ˣ$���۔ ���r��-��z}�-�b�$���xbrn�"�}�P���v)I�SƵv�Fjѳ�ɏY����4g�
�t���y� �36��Z~w;��߀y�&�ئ���l{�(�a4З���ct�{�-C��Bu�8)��b�!�dEO�^'�fD"�xB�"n���Kj��-@CQ&�,��&ȕ�A	��2�-rnY��:������[�@�CIȸ��e�_Hp[�Jv��>�%��E�-��Y�5�ܰ_�D9z�[0����mG2������˗{��f�	<��A� ��+���K36T?7␫8浮�*V�m�u�S=����J|A3�!�G�Ķd��V�J Y�E�e\���U�KS�|]�4k��c�y�A&�ګ�h�[��<���-{o���j��E���D��&p����T�H&�Y�p�K�ΫQp�Sq�wّ����7��KX��X�=(
����W,��#�ߧ xO����ּ	��)L��;&����|�\�`CT�C#f��Ր"?`Q����x4�a[���v��H�"l�_74���	,qJ�����@���gr6|���|H.I�$��Д�d���$��q�s�][��-J^��UZ�zaI�)�[.�
ꐯd�eNFl;�|�qr.7��Ƕ!��aj[[�}m�S{�֟�H��4�7 �ӿ
uN���4��m����ZU�
$���L-�ªOA�	;�>�]��1]�?|hNw�Q��۩i��fp|�J�|X�a�#������'aN�ۦ��������鸵�s��Ml�7&�Du;�n��7L��~��
�G7�|�H�[��?t�`�N�=H��Ǒ����r�lFkC�s�U���*ғ���U���J��@��=��o�ڊ>)3O�{�U.Ziu=!Q����	�Q�2�ѝ��-�����%a8W���
���S�wv�PD�vk�������^aH\�c/� �GɌ6j��r+0>�ؠ��%��?ߵ����p�
Ļ�H%��fN���[����r��k=��C(
-D��eG�&T�\�}n���/ܡ�aUʐ�aE�޶i���+�$�s�d��g�6U�摇$�f��m��Q;/�]w��d˜&�v�I�P؛�87B4�}]<����}�p�.�n$����ϲdJ�����U���H�鲨aת�`6@����y
k3S�u�'��'��`���gQ������.+��O1�(D![>3%�=��o5�Ia�$�����<US��KT������u��l�c/���Q'����m���۷�Xt�T�5ǆ�;`h���&�,�
߾�a�'Iz^nAK�}��u����g��3f)���g&���-?��-D:�fY��z�D�,<�8'6�^neJ�F�>ν�A�!���\���Fe��Q�a�9DR=�DG�	�&��o���̔�Y�q�n�L��^�B���jA<҄���#hc�,���9,���
�M:��˲	�5$|�8#�n��F(`5gq����|��:����N�i����ҙ���PȜ���k����OБ �P'Ey{��z*g�j�2�^�]����4�28�xfgh.L�/;��ڧ1
D��|v���c�^�/���ư�wy���,���n�nk����y^�F:�b�"�CI�[2�X�5h���o�ή���r�'����ͥJ��7��<��g�p�-T���f3��^Ͷ.qiD}��*�����kIJsO�;��C��_�j:[���[?��B\GS�=e�*$�dn�u�ƺ���A/1\������ry0�1~�C��,�'ކ#+�=���*~���I���S��
,
��ŚN������5�t��R��vy��G�:����rHc�h[�X��'��՞��9����sK���C��*����^�M>��V�~�_�A�>R���[�
)x�T:ns$��i�~�!Lկm� �K��w6�ڮ�D�9�3�0��6���\L��I����S����Z6T����1}�zO)�;�6Xlh��B���ݠ�v`�<�iqr*N�+~�g`�ƉVx��f�e��y)�]Q3����'[�U��0�F�͵�6�W?=ۭ(4��b���d�@�"�^�`<��?�DC�p=n
�*]�:1ϹU����e릺]��G]���,�1�<�T���~E��/?54PAN�=��D�,j),Lr#v!���H��"*R������2Kg�|�	�m��(̻�ϊ7���B�}|�LM����3_j�ac��^�b��2�=}� ��(=;�q�^���~*��g��)�!���3\Ѥ�~������7Ć����|�o_�n�F^,6co"�����A�~�@���8�]�5������A��.�G)���]m��& �B�j�e���|d�غ�^Tg:[ݒ���(�^����������b=��Қ���F���9�;�Ł�\��l����N<#�zg�� �O1�2~ˣ ��꣭��А#�Q�n�빁�H	n�`�:�APQ�Y����{�ZP����C0�0���z�c��[F;�ҰMҪl}^�Y2�iйN�BZ�,���?N	݂�n,��iX���f0h|��֐�,s)���nw���]�Q�I,�5��� m��E��5 �8�c,%�����Qh�R�/!
�$��k}�,����'G���=U�[��#z��ff���^/�]�Œ�S��<��̺s�3�>6�=f��{C�f���V��YQ?~�T���c�k����Im1ip0
�W]'ב��y�P��͛/�*���]��D��41_s�)�*�V��I8(qҠ�E��Nb���1A �v�Ķ_�� 6���@���ZN{).) h� ���Fυhdp�����iۑ�Z@�<�&��q���Y�NC����[�=�x�bMg�.r�K�B_`��U���u{ec?��Q��Eο�EoZe����1��!3Rb
��(���W��5�#�������*�S� ��,�p��4���6��_������V/��ۨeB��3w����0�-Ra�d������h33Z E���~T/y���S(���"A��+����u!��?D�k�5�$���c�N���н����s�-�ص�e:���S�-{�M��������)����\��5�N�g�̋�[�0>�ƙxg��ff亱��9�)�C��@%&"�!�nXZ_�&7"�
���d]�p��j�)?ʗ��������_�NEe�ǱN��d��y�+1��e}}v��mҶtӂ�b)��\�b�/c�*1�w��Ы{�8��4m7f���$y&߃��m�W,3L p�d�/�G�m��F�@�����
��@�Fh�mf=kLrZ���ZfXT �ӛ�e[��[.x��h2Y����**z�����{�ꈛ�M���w�9`��o쪆�,`ypn*� y�C|������P#���6V�j����4	Rע��(���.���t�t>�p-T��z�H�载ZP��v�ƘP;�5lt�l�y�yGe�ێv%��	H����<�jǨȭ�aFT�E[���w��k�#� }��Fg����V�R�Os�ؿ�y	I[G'���WeP��Iȭ���f�@7N���'e����]�:h+�Ú��v�������TLJ�D�D�r�dI��d�ڪ����m���kw��@�����:0k"lI5��z�~��"�v�Rv� ��|mɸ尣��kE�p���w�%@erZ���,��/>�д��'��X����\�����|�ai=��+��Y�k6~�U��h���a��,�C��0%���ڴ߈O���ӭ���+@8�����[_P����C�nx���x�[3�a?Ҟu!%1yU@빞��r��=%ju�X!��5\��{�*�{w+��<i*)�<�վ�j����7��)M�����:�@��cv~P����z����Y:WU�ȱ��x�P��LS��G��.|J��N7�����-O�Z�����vN&K���������1۟����ɼcX��W�5��O9�_� v-��賚���a�}�I�3D)�%����7@l�� ���j��P�FĲ��/�O���&P�g'�M���;�=6��t�9]��>��$��2�%�ĩ��gea}m_����x��P�����S�uW.��;��%��h{ꮏ�[1N���m�܌8�&�����*�Z���٨�jqs�V>�4�4���Wi�F	x%E ��@�֓.�=|_AuK�Jg����R`�l$fᥴ1_�VY#�v����E�옸�q,�������Tj����W��)�z�ͳi���ZÉǑk���/xāt��0*�W�t�%� ��3�-
(X}pc༱��������M���֫EL�[-��
!��-F�&������h��D��(74�fCSn��ǝ� �5Ԙ����fB��x}� J>��!i�@��9��}�k�ʿ�a�K�Tb���j�{�n�|]�"���u*۰�A�I��-�C�+���⺳D)T�I����ٕ+S�F����+rd��/�w��K���ͼ:����0�(kA."��yI]�Q����ֆ��{�����3��񹐖	��dq��ի�]��+d��+o>��\�ݶ潒�{"��qt�|�T��@<`���ْ
�ZC���G��u!qj�������'H�����s�`�F���������"a�_�R��S:��֪ؿ�<*��R"�l��GYPR�|4a�t�~D����H��K	�N��,�������}W�;�B�����y�@�A�:$�
�j����4@�'�4�$G�J^�$p��8:=FR��@Ba�22�]9T�V⨀/�ĸ�-s����YNn����o��(��u��թ�\;��(�<��
o����{��!��t��o>��z��	}�R�T��_1�e?Ŀ{c�q�E
<ݼ��0�2�c�� 7��1|�)�m��.?��~�TH!�I�z���9URe���᭐�z�{iѸ�e]�DxG+ľTǈ
/�B���FpK(i"H'$M�鴏���k�[r���:LU(c<���?S���$�>���kK�Ne��r�1�
����I�b�0�߼�L��ȟ+ �������q�7��Ufs:�F!��y<h^�bR	�M�,��&����$ղꔩD�������̐+���(��'��~����x:��&ϝ��!�I��cU�B����;������D�|�:�&I�
S��,�\�[.G5�����li��2���<��0`Ǭ�����+��]�^��*�eL�ċ=Ō�Î	�R��gZl'>�W�^]m�>�a
�(7��n��oa��aC��q���hEvD���;a?۹I �f��2!ti��ej�A����e��
2������_[��kAz�dw�"H����6lݕEp� �N&���d��� ����$���������/��Xdk{��eO>�[����@������s�c�(���4���oY��J��U���ѹ�Z*Of������	�[Yu�.����߽y��D�7�Z��	�V9��=�3aR�	Yi>�J�(z�G�a*1�Yo{e���)��A!#ӥ�,ｸ����W᯶ ����ʶ�Nl�a�b��D����?{Q0M�֬����X���o>�x_m�q��R&4[H3���#H����߰r��ȅ&�q��:֣-�l����mpjU�^�u}]o53�T?4g�@�
!��QOP�1w���|��k��6�5R�6��.L%� ��'�\
����L͊J-�y)�C��pk��3cɞ��iǒ���q��z]Fsߵ��W0D8����pW�݉}2,
ݴ��0ê�N�Al��(�6za��s�ԭX�u9*D����m ��U榄X_���>*:��9�U��/IA��cu����`���=�m�Z��׆�#�<�e��cԡ&��k�Cs�զ��Lb�wot�����A���p&K�s���;�>��q\ke[��E
q7������}s��I���5l�:��~��`;ќU�����?ݖ3���)ӣ�6��`�������>XK�l�;G��s+�Y�16�����[x��c�{����/�X��!�
�Aݛ5]��n{�Y������o�4ڒ�eHWfO��mɄ���0OÕ8t: n��He�@oy4t/���8B㵸���s@��s<T1��.QM�Kʱv�t ��(�W݂6�0���}:B��'�"�������ޅ��a�,�'Bh�C�!wFZs|�Y!ޅ3h�݂����&�����R}��Q·��5�D�|��MpG	��K�)�vڅ��v��C3q�/!3�.�}�t�8t��ܲ+�ϻ��`a���Я���gxtU��m/4K�Y��;Vf�I�X>Uv�>m{�����$20I�rڹm,�cM�P���c���b(�'�/�iP��&,�$y&)`Ӂ�7�e�X���:�{,nm��f��Dt�ql!�If�B%�����>υ�ox�>QHߐO�-�i��T��^U7�����@�W�
?@�& Phy���6�*]�21��[_Ȇ���S���(Xbp���ӽ1�8�&T����b�t�J�5%��B��5�E����"�#��Z䓎��m:�_ۆ� s`�J2pD+�T���C��#]reny�D����#�r�B�)�!ň}��mꓕ+
�S���f�uZ��5��|Ѱ�/{ǯ�Y���p���]�.hҨ���ȋ���#�K���A��g�CjwL�q���_]�5V�4�a�47��ԇC�?ߞ��t__s������� �"� ��򺚁�GO=�(�|[Q���O.X�gef.�vD�r���{V�K�m�5&�ݑ�e'����Z�D ��" �~� yPK�;����������s�m!�d���'C���9�
a6 b�ȇ���;���t�?�2�fmp���4�k"~�	�C'�(Xj�N�T2�Q5�2Z�5�ٷ<04($�b���Q�H:l�UA*b�;�~zu	��E�j��J�X֏w�Q�"��cL}T����PR�dp ���%j٪sR�'�����c���O��}	�������������- ��1#��M7*ܘr�}�Z+c�?���8�h���������S�+����N��şMY%ܡ-UK51�����c(�VD�0���;�;� I(�S��j�4�I���a�^�$49���9�F��Uۣ�S�+KUQ��@޳��xpg�*@�����~��e3P)�DG��Ӝ��Ⱥf�#:4����S��p�@�*��/�كn0wq�(vL$q��Ù�������|N�4��}F�y)J���<c�=�rz������@�{�΁6���$pz:/w����R��-̩��'�MF�E�����}T�{׼��E���v����f�;�^�mz'R��F�:����~G,�����5�;Cr�rM��GE��#�f�{��v�>�+T�������\��̵4b��U�3�x�޻�� Q�k�!��*f�6a0��(i��3M������tǽ)�G��hz^p��-����7�7v��=��:H
[P���Z݄w.I��R������V�܎wY�UFEr��Wz��m�x�(F��� ���L�?�C���s��J���v�B:�� �!G X�tM"@0c�	G8����i���t�s2~;��j]��d�(I���ll1�1~'�$�g-ǐ��{�$<��ꟳE ��
�<I�^��jܹ�+�(����x2)���42�O=K�3CԨt
��P����EK�n[O�]��b�WM[@Ѧs�F��U]yԒ*��z���WdС`V�vy�lǚ:��L�����BBnR�8�(�g�6�A���r�;J�[��備�2��v�ĎA.5�A�����.�P�|���$�J*jIb�*HT8��EܗI�|�_��o˂@�hb����E�`(���B���Ҷ�gbX����/+?�ND���_��,5�2��	�VT��$�Xqr��JNX~�>W5�v��0m������]�SW�a�Ԅ-N�ٞ�&?A�LgD�/���*6�%��/�rZ�8il`��vŹ��p��l`;3�޴�j�b����T(�G}�����K�ZԂ`LI��Ye/E򷚮E�M�
A��oN��Qt�m�{٥$�����78�VO�!�vLL��ҟ9��y?6
����!bDo�8hVo��f�fd�[�<�'Qi���M3`�*�A�'L��@�U�J��l���p�����k/����k���k�~�Iy�mf��:.�b��*I�e��A��C��,�L�+�!�$`Z3����DN�H��jw(V� �!�5�>\r٥L��
$(�^�f��)�+q�!�־W���d"��8�:?kF#?F�`c�-e�yI�$g{1=�]�KҬA�y�W兩)VC�8��i"td�R5��C�[4��H0w��)	�[6I�a�ZH,��i�9������_քT�Vb�/ B�&9� �����g�#�G��!����A��st��Z�q<�7��C�0O)��/���g�)��~�'�ˊbN������P3hu��m#�v���P�,�"�g�%I(��\���Q�����.H3��*-��'��P�  ��gjEkdE�L����K2��H��}�e]a��@�}��)Qz�LYg��`�C���+�yC[JJ#��#o��q!�3�
��&ݺ�}~�	�a�l���}Վ�ΎS(�+C���T9rF��i�u�������Ѵf����P	��6.�iAe l�E����/����he+�SV�
1���w
���+| �q-��Ym!i���*���ƀ�벦mw���)K�D:��B*F��-<"b��U��e�.8�\ ����(w��鏨�
T�I��>�pCz��T�,z/�,��Uz�D{� `mS/�x��%���u��d���M&`=���dl���DM��s��fe5��0����٪#���(�>�K`^5o��$��f=�z���e�� ���>��6��"b1}�7�k��#�cf��Z���CS!K��N��ax�uj�������mݶX�=h{��e�vԂ�oh*�:H�o����w�B�nT��5��Ȼ��Ho�&�ǅ��츀�������v���M�,}Ȝ,�ь�?�����\'���-�����0x�5'��R%�e@'N�/�W+�u��k�ӡ���)E"�V����9�j�A�ED�3��'4F5�`��;o�4�=��I�3���@;�[�8��ƫl�\h��Ӷ��J����=
q�]���!���~P����~���L�l�@���5�|�?�'��YK�?�$�_7_)zb�,X��ն_����4�7��;O�3�{9��:�q�U��`,!�W�����r:�$��!����_��O����l9��6�B;۟�b�����9يʄГR���{��G���d�����d3e���-�ڑW`�%�]�tI0��S6�*�I��!<��ϯaL��TAn1$Õ��??O�3�CnV(�� R��͎ۭ���evj>|Tޡ�B��u��B"I�� ����O��H;n�ɕ��_-Xv�1�	q3���?.���N/��{H�&���Sn-�<^R���%d��p�X�&\"M��eE�wp�p_�! Pe��:2��u�m��:E����U(8��(�x<� U?���q��&
���X� ��\����RY�^W]B<E'�� !&��"M��Z����F	(�m�Ku/�_Y_�(�'�^�*��IV�N��MH=���2���
�g��ՌY���Ђ�k���U�����bB�u��jXb�j���1���H��4LXۻ�Un�ʰ]�?�+�W�d��F!�s0J֤91�O���I���:~N%�	���yn�E(����FP~����8�3)�Or�!�:�s��6�p=��IO�t�ftR�ql�ǲTI%߰2�uŊ�,��P�"4�����w�D���������	��j�m�/k�sF^�}ʹ)�_Pn46�p�f`tR
?�}ZBZ*=����u J�"��F� �Lo>z։^��3����FD;�.��!QL��_�%
B�5����{��120�c��R�����V�� UKB*c�1��\׊�P��;51*kO*��OeJ����Q�mK!��'A���-�����:/�� �����O㜵���Ep2GMk(�$s�Z\C��';�촒�ӿ�X�b�v����	�&
��h��P\�lHq����α�i8�2��31y:��QQه�ގ��B<y��)�ڿ�:7���:����ù6V �*�B(nu%}�]B��p�0eKk�>֍W.�o���V�EQ��n�R�e.��I��`��Ì�GW��7&�ET�}��5?Iy*�y�(�|�+�$�$�'��R�W &�?���V8ef���ʗ��3�yNc�;��g%)ԖT0ۚ	�n%�{�����pGV��Q��g,�p6��g�J���
*d ��� �)3�`k�TKZ�'�#ln��8 t	LF Q���~��`I���U��Ph���5X�K���ba�`"�=X5Ѳ�Y�д?z�wI�U�
���n��}J�t�����Ԗ&A�Q^g�9e�d�ҿF�B1��.l,NIRA^XY�9`_Q�5*�9*W"��iw��_�>�FO��ħ�ԣyd4.
@�k	��E�Sdn�~:��ܲ��b�������Η����wr��<�������L`m<ND�Rə��YI.�3ѿ�?6����?C<��3�x��T%弊��>�똟��@Vp;hvo��ܦ�e,��(�:J6/�N�+,�mG�#n��̠���T�u�������׬��nDj��If�
��&����hDr?��B�v��9��W �����m#���o+V;u*����		&6�*`衖��ٓUy��.��:�۴��+g�P͛�;��9�,���-�
��@{I%k�՝lw�&u4�R;"�`g�A��mG�V�{AA7��iL��!R㋓�h�Bg˱�\2�k��q�n�8)�o�Q�37 u*߼��
�����??󵃐��O��Fəi�lh}�����7}N�LȰ��Tb��K��*ld�1�jF�����c E-1��]L�+�E��p��(nl�5srR, G@�0D��)�ϕ@��n1^l?šQj�6�}�v@	�M̈/v��;"DVg~0M|��LN�D_%c�(��\���n�t%��w|��6_��#{O�XR�W8�Cc~Ԫ.Z���{��J3��A�I���Tv7��.�+ld<�o���N�/�x}/��.#D|�V�p�y(JH�؀@��W��B�D��J��R��8�E4�q`fm#F�4Y�����3�L�$C�>q�"�
��UG)
���:tXBoP�ЃV4�U�'���p���$�A�,L��������A�{�5ϱ��5JP9�*�:FfD��@&`\�i��IMh�@Al~�
�q����A��Bu�X>S&��#/�M��^I��6�u����)ْ�js��.��3Q+HVkq�x,H��UK)��$u���?��I�X��ɱed��,��2�K�<zv�:��5�~֑JM�P{�%C���T̺!�;�����$]��^z6�|@. W�^��=��i�RB�7.}��_��!&�=�A�]V���V�Ȏ�^9��aǖ�%�k-�T���O����B�����k`_�����F��*>&�0HW��%4����+�)߀��d�p�ԁ��z�n�w%�~+[�B�_�=T/�˻zd�1X���u���m��嶝���?���.�+�9�g����[5�����O�rt�ܳ��br��҅5�@�IA�����^�r�?��h�'���Xlxc�ă4���� ����oH�Mu����K"2��t�U��M�T��1�U"����ɧ�%q�nܛ�t�����J��c�q�nH�n�P�<`��lR;�^� ��ƿ�����]�B���D������?3�A�ؤ���*V�Y��J_�ԃA��y���@T{��)||N�R�Ǩ����|��Vc��9�4W���a��x��J�*]f������C�,��뵤rX��ZR��!>�K�ǃL&�����Rk*JL�x*��C"R�׺J��Sw�]̢�`��T�5$����{�p�&�T��ɋ��)7���e�{"��&4��f�����d��DJoqe�2iT)�[��ݒ��e�wn��錾�h�����Ka�����Ю��k�����3�}������yѷl?oe�`��6��p�d׀wU�o;��x�Ƞz��~����(EP�X����ø+�&p:�����NO��.��zl��U=������N>����(��7ԝ��s���.������t�heC��G�q�[�<�V0Ŋ�ou �/���@���d����͹D w�:�;�ÈSQeJ ���	w�w["�U�*�JwM��e��m�^�������<��K��!��9��S��ve��m<\6�P�-1�	w�`ʅuw��jf�9����A��K>a�:N����-w��.�18����aZ��Z��{`�ے��>6Ն�<8���
��Ҡ;\��a��hG0�#�{�A�8@� 丄�G�O���~�K�Od�Ӓ�u�� 	bS���l��8V^/��ހ����q(J]K���~H)ޢ�[���?S��ڋ��_L3����/u���w͢6��@���ٴO�hk6O ��C]d��vf�(�i�3 �,�2YH'w?F�	/�8��o�<�Fۡ%��@V��a��W�Z0�y�!ˍ����"7�A���#��n�ղ��8J�Hp[�h��f�����}2���>�Ly:��` ���E��}K����}1Xe�lvj�wϛ�Vn�� ������	���8D��Za����6^ ��-����ߛ�E�F��N+�v�\���$fl���GK�0n��jo/c���3\3�5�|@$&{=�W�jԋ��9tQ���t����-�\&he��f'1e��Y��;��g��ܬ���/t�6��P�Hu�=����R���7p��3y��;��#�sU.��]R ?��47&�8q���8�{Ϡ����-Z6��O�e��ѥ�+�P�D�]UW�`B�9VSFg�j)�(zݙc4��<��w�j	��D����;D�$�ƚ��GM������Fo�`${v*+6'�c�j��h}���h���0��xH���.�����?bd>��k��M�l�do��[�aV�m�gD[=4�u�jL��D��ߡf�:��b�>�̑�+V�NQ�3����<�UФ���VM�{�и�NpLt�T�`E��A��[ª�x�Qtݾ��лX1П{X�wi�͍�9�m��s�1��)�&eLH�P�#1^*G�|��8��}��C�>���k��<>��9kHa�Z�,��w�[�4�tԘ�q�e*~r�`]	���i����y�D��'��� '�P���HA.R��E��ӶÂ��f�L2���jU���41�ff>�ٚ.����-�6�e�H�fu�{���$L3�D�����?E��c�Q��dr����=ܘ����+�p<��b��M�1���Q��9<:g.�E�5�u(�����Jhd�g:���]�Dv�f�^�4��u6�h_��.��� �ݾ�"B�#��SQE������{�7b�����������ސ�
�]v��,�P�����1�kO"k�9tuf���|��gS<?�dSx�����z��m�����/Y;qȖ�%�bd��Gk)x,��f��o�;�}��R�9EnP~�6h)1�P���L���w)���_��b�S��<
T?��x�gE�%�	B.F��B�yͳ�o���c�'�nbBOy�>q��,�h�����=i? W����BF�؟О
��'V
b]_L�	��%�BF��P��Z�\4� �FWxl�W	F�Sh�Ik��1�����q�>�MG	}�/}�����{P8�_vMm�b-Y9�C��%���v!�ׅhO)H�}�(ؼ�7u��윦������ ���/`6/�h,扑nY��[,���Xl/D��x�؈�tJ柤��p�Bq&(�B��Π���$�y�D-~:�i�\r�k��y����K�ψ��2�`"*��S��s�)�ϯ�JI�$��� �<��zh ��\�B����UT��rj����NB�C6W:��y�xB��~:�3�l+�o� ����)H����#�;�A����ӛn���ϡ���t�UFS�-���@�v?V���:�Nx���_
�����>��O�a�M�r�TL����`MO���C��^��ZF�^?Q��rl���|������m��"G!r"�s���q&J�����	��tf3Yj��ٮ*>r�c�#�.w/��2���L�j�U��I�e�:JF �PᐔO���&	�H�,K���k
d������� iu�@a_��R(�ȭ ������R����_p�օr�������B����#�-�!����؉_W1��y	��9S�p�m���˛�p��h�r˴`+M�)�c|��ox��+�[x�,~�F:տ�fC���8t�����_�}�!C+�fb[.����!Lr��8:%�.p_��~���5.&:ڊ��N�oZ�g����lh��c����|5co�.ro�K�!�ʊ��R֨6<hj@f��hQ`{.�V9��Pq�������&t�23�}��*�F��f�rf/���ğ���;6s���f��G��v�8�~��(�(�Gl��$r��d@�/�lc��	�%B�}��	4N�^:fo��KA7G��~n�l#�,�	�DҟG����=�+ �'�P �ҩ���uj5�!���2FaB���y(�R5ٗL��)��G�F�3N�۰��f���V ����\ߙc��`�6��(]ſ�f�W��>�Ω��#��B7ؐF�����rb��qBz��	D��������E�T�\�0�S�c��`�3���򋟄 �C)���>�J��.5RىՁ[�b�7r5���Zxw&�t�T���y0rs�w/���a�0�_�( &��7$V7s��gB��tT���Sa_��|�ت7C)oJ�A��N� ?�Xsɡ��[7h˄�ѻ/`s��h��͉CC-W��)��#/�	w�KL.Ἁ��,�}rd�mW�<M�pY��bo�N�S;����s��J�Z*�!�XƓ`��=�nc��zȳ�m`�m���l��~�X���m�(F�g�09�����q|�xD�ˊԸ!Uؾ�;���m�y��<�}�@ZE�,m�Tn�ٝw�
>�)�3|��?C��m-*�����-z㩢\�)D��a��nnn���  ��&1�rn�f��!�wv�[-h\ �9�!�f����T��0���$O�TX"<�'^qs��G[�H2boZ/Ztf��|`DC��jZсF<B}*eHs�o`<��A^qN���H�G��t"ӿ�E� �d�i�*|�4"џ�<�tߘ̤�4zPy�4��a�a�K�f_5b�M��l[۲�](H�����v�^@=sg򎢘�^N�x��Cct
�,g+��K�8di� {`��Q�jP��}A�\�7���=�X�?h%��3 ,0g���⬸=7a,��=�N̩�3
FDix�a��`@��{�0K�ࡆ���I�;->�7��l���gA�P
-n&���!�h��Js��+/�xۮ�F����a�<�$�<˓P��1)��v��&�����-�CH�36)Gh��ZF�w��b������V�"��}j���n{�4������@yZOJ8~��R/������t�9X��K(V}�L���'��9Kj��C1��`?��rU0/��{s�neW��*��F�`�B� �,���O�a��܅�e����3lى�<?�nL���#y�w���y���5`6J���hx20*,�W���,�lé6թ��������~a���IHm��Dy�f�..-� �XI:?R���J]��o ���
�����x��P�]��1����Rl�f58W9��掬J!���
��wf �D{�ϥcU��<{�L��l��W#F��9׎Z�t^Uf�^ê��vyUNG������J6�?�1{JOj+|8��`Y��w��*�_���5�X�`�<�mih�f].^;�<
�����T �V�4ω�����N3��ļ$}\��x��͹���f��b4p�u���H�-�m*�����J X�ٍyZ�������U�;T��	�1i�>���/,��:7� K��$N��a����c����v�l_h6}M���_|�[	�i@��2Q�����m!2�S3�QJ��B9BYK�n�7����(�R��W��G��o�y��G"
�0�sb>Jx2:,�	nեɇ8#�3��� ����1<�_��8�Q�:;Y�l��1
Ex)�c��G��GDK+��z��j���tv)X#�=��|�c�Y��C���$���Ŝ���9`u-�?�����l ;[VB�ۤ���{�r�G����s�#d�K���Izn&#c�>.,NO�R����Q��g������$��k�<Wґ$���I /4�љn_����sI���Io�a�2[OĦ�a+�P�����%��Ӧ���x��x�"�"���PĜ��� ����MUP�=�ʣp�"����+���qu���蒁A�(\Y��D�pX{D�C��?(RL��*�r�#ߣ�eo� ޅ0��4d����Q;������:����B���=r7ȧ��9���I�u#��r"Q!⥫tB�D��`<
"0�E���J�l�H�mr1:m5��-Jp��?���PH�M���󍕼s�PU��i����?l�2�P�4p!����85G�n��E<��au���3�ea2c,���h	�s}RdIOf�}[�ʣ�K��RP\e�<魌����Ө���,H?#�~oj��>X��J����5����}Q�ӛ�+v��޽=��m�̉ӹ�²��ӱB�Q/@I@y�L`̑�e��qгі��N�u��gQa�3���+p�u�����|� X�L�����LN-{��=���]O��_U+C����?i�<)��R��k��򞍧A�i�H�s+	��Q�V�){,-R���$����=�\���9 �5�-�r��b���C��#ي�--4i�����_Q0
h����}���۬"�|w��c�]�,>lJ0MEg��~^��?��0�D�!1<˽X܆�_�XR=�#�6K�}H_,?�m��TV鿰 �%��gQ��N�aUnEe!'�u�h؆L�S�o�|<0�	^��V���<U����Z7�N��f����O��ޏ��x$8����rj�P����mݹ��L{��n9���p\4��%+y/��m�;��u���1h�+uQؤ��[B3��-�`d��(Z�Rߏr��֧M�Qk�B���&F+k+>�GHw+�t�h��:�ݏ��z5�o�v�@��C)M7�lg�=H&����sԁ�F�M�[@�7����Q���4]�$�y��ST;,��e�P�D�����'���S�,�Gu���S���3��Hr� ��bX�Ƀ��%������zx�!�Ř�M����+����+n�j1Z��*�ވ�{w|4,��p@Q;���M��Qu�xRP�d�b��T�(%iT��Q�[-�T���Ç|s��	��X/�m��O�v�	��;w�TX�t E �W�g$k�������4����!��g���:������d�z��� zBŐ\��K*K���5l�C�}�jH���B�X猁i9�~S�	#c ڧ��8��w��-OS�_�E�8��Ӎ��0�΋��9yQqMc{
ղ�]�+K���tH�콗b�ʦβ{a=�� �Dc� A}̯ng�Nרw尌�P�c�+�>����_��'����*�we�{����a�V��<�~P�M{��ү�y�v:��9�0���j���sq�7�f�E �	�e�H�3��]���&�����)��F�%��S-�q@\U�+�=6h�͚O+��Z����g�KŻr�	�v���d)�:���� �H�v���
��uJTw��c�]�ZeW�Ñ倩�9��A����?�bG���,�����ትب=h��,���s����b�k��Ǒ�g��>��d�Zգf�V8�n/-��,��Y��g��?��5�e�̐kL�Ä&<�Ugd�J0)�f��5���%����'�"�Z]���\���?�b׊G���_�Ӎ�S�W���$6Yz� ��Q�g��g##��7/+߹�O�y���Λ�c�%���o�4ژ���i�kgM��L�I4L�? =v�@�LwNu��I���R�!jX+~I��*�|or(<�`8q��ݭ�p4@�m��/a�Gy�b��u��7U�9��x*;,�$��!�&d�m$����K~�w��Ka�'���/�U����Dn�A�EW4�3��j���A��R�8�Q��/�&�5@h4����ϙ�5��t�y�|T���<N���H��u��h��Y�q�C�����Y}D�Z�9���U=Y���}�7À�W�vz�CΙ_O�!d(���l�a���!�aꬊJp,B�BE(6" ���R[�R��N�3�9-n��V��F;����X:�}Di�a��5�8�&��N�bS��#{�n�衸v����d��K:��j�ڂ�q�>iV�f�9o��/�
�6]�Y�F]���,�� �w,�)�㄁��2��y�w'������$�������&���|8�+��-�P!Y�G[��4t��(6���>����~�u�m�"^�K-i�����8�����%���ތM�>�;s'`������V�r.w�O��-(.�6k���p%(�L�8�k`;ڸ�� Q������.�?�o����kFkX��Z�x�c>����^H�n��K8��i��L�g�����UQö�.��-�4Wj����"��?���}=jSy`p�P�����:6F��n��F�xD���2*.H������U���7��H��{�"ܢ�l������3g�/^f�HaN�L)�r�.�/��� :0|�c݅��0�Z�zcz����Op}ES.X����W����i��+� @�������U��sN\��0Q�DHV�3c�C޳�2xW#lC"=��z˾����9 e`q�Q��Hi�JE��|н��%�h��%�goZyȿ��u	ԝPrǀ�2���
����ٝo��T*�R|4�T���X�ahhX ��� ���I���!'���s>�*<������hA�-:ϷPV!�xX�`���W9��0���2��U)���7�ؓd|�+�9���V�._�>^z%Jm�w�>1�16q�Y���3�;@���rM��5N�F#���tr��:30[������Gq����KBiy���m}-��f�B�_�bc(�ؽ�1��Ԇ�e�{�<P�����0뿴�R	�u�}��w&ȨB�,��)�uO͖���0�����ՠD���a�h�#�.6���P���t���"]r,�r�dP��i����Q�f�}ܜ >'��W��2��e��Kr��]t�
Z�H������?���}��s����
39� �u�� gg��̎���隹t˝Ni��s�)_�]�Qr�T�J����s5�]@V��'�� �|�1q��%��sT���?.Y+e7�����&e4$�X� ��������剙1@H����Uaӵ�9.ق��-�F�i@d�\����!D��y>58T��ᨿ5���.司��VQE5�!OM;��e��惊����Xt����.`u5�4nu��R��)����"5mO�(K�P���"�f��(D�KT�I�#z1FM_^&�$��uF���v�*$?p��乮�ߚ?�M>q1����=b=���y\h�xa��0��o�5��IQ8�6.[�)��,<H�-������|c�ȣF�՞�S�?x��� �/������޴R��D%v_"1��X����H����8Xj R�ټ�G�^�!BP�J�o1�f���[�N 5�b���r^`���1y�zu~�9�}�阾jP���FY `������<�VCz`���L<nd�O�L��I>R	 [���U��{���o:&���5������������e�c)�<�a�Q������\�຋���ۭ�����k���""�7f�qD�e�C���Q$���3R���� 4�����Y�\�|�$#�J�Lr��[�s�`�ժ9-�م�;˾��at�n3�m�o�ZɉB(_+���q�LR����������YrP�Z�z������Q��y�/b=2�D2��(q�c9�}̕�X��(�X(���-��FSRZ��l��I�D�`L/^WV1@�x�f�� �Φ�k�i/���\��Aܣ�`$Ɉ�@2����	؞�G��/�r��,Q�K,5�����ͮ��R�FjEΨ�\d/�c��E%���)�h���o��/��h4�Ų-��r>9�֋�[E�ڽ�}�˶'ˉ�����C[L�{}f��{r����?:$.F};����װw����l#�����4F(����; ����j�U�*G�o��X�#U]s� w��,�5.}:#9dVn��sI%NZ�������2s�4���`	A�C@ʷdW���+���@�ey����sς#y�	�5yg�m��G��7H��c	ز�YU@�*,IO���NQȮ�q�[�]ËԪh�2��n ��2%A��4���FbJ�D{�>��O��X,��"��4���mK�t��@ ek���9͌y�@%��%�0�{y*.�tUq�z(����I���ȭ��=S���*4�`��Y.Ӕ�ԁ��=u����WO�oar<�k����@��*��W�۸B����!�`�c�S��ĔZ%M�ʄj�F	����ߕo-�9�� �tʤ�E�+�r�Z�Jb[ߜ�*���6�nw��S^97�(���T���M�$�!�����6�^B�l~�x��ym"vꉽjV�ɯ����a|�
��ħGɉ�4O�I�'LP��G ���!e̡�[ѹ�i=q���Π�n��~�'b�OO<&*({=��ֹu*КWl�?K�'F�X#A�!��R|!���@s"êڥ�`� ��N%�3�������9_��^X�bbJ�0G:p5������#e�����2�d��FZ2q���{p�yc�?��b�9��<�q8nݍ��t2 $R:��� ���^!u�������,���"��qے�5`
T�����
�~�D�5��Z�U�u|Y���w �y6_BV��e�I��[CՉ-�|5"��)�����y�}�-Q;�7��o��.�1�ݑ���"������(�����g��?}ِ���)��_��⒂E��Σq���KZM�	�q����~)�>p�l\h�_����$\�hN����'��8�=���.I3N�����2˿��i;-!q�giPXB7�P�������)H��԰����S/H�
�$?����(q�\Vn�!��&kU��y��l�c���:ط�:���"IzG�\%����joT���C#����ܱN1ef�T!Q���
~��Q$�uM��S���0�̗���&�<ū�����}dRq����)�
���Wbd������oLG�T��hpe�F���7�,����U����F%U�p������<6y�zvHr90F�}5Ʒ#|�N+]&�NOM�����=�0<U*����2D����w���$˽����:�	o���j�Gbx����A&��6z����K���%�R�������wY�{��ާ����=)��������M�K�A{�1�f)��
$�زZ&�(l���ͥ�`��4{c^~^��c� �ۜIѯ*�M��~ �΢'yl'�_�_���#��m)�,��![��qIٯUSHOdԋ�R�8;�,�/U>`j~�ffũ�2]��IH����g�T���_�̖�^tp��{�����m���?�ɉ>.q �5��YJ}P�>���Z��e(kʩ�o<���-�������A\�S�c��:�˶�y�y(^ŧM�z�:5�����p��� Q��
[ P�F�[F1?zS��+)�f>�>oY�Z;<�ihacd0$z4S��o�oC��f�����$��z��q�/�\�]�@-Yo��y�OC�	rIɠAT��j$��'�Q�Bl��-Ȳ�7��<��sÅ���֖��c3CYb�#t� %*n�bSOz��-v�xR�9rb`6t�!4��6I��:��ֿƲ٦,�a����!'�ݗ+�Ģ33���=���s���ӥ� 7��0��_��c����qG��g�s�¯��n�.���pe��E/eTm�P��dKx#��z���;���V�_��B6fjQ�r��5B�N �A��Iu���`��_�,%��\p��m�;�u\v8~6�q?��l	)k��!'j�uU��e'<#ڪF7y�~#��j� �Ďw���� ��ܠ�o���	��FY>cf����e��u��u�b��ES3�#��d��������L=?M�� c�~�Q��6��,�l�Cf}@ˢBg"pf�5Ѷ����$*7��ڇ�3�8;%�[s�ZE�(j����k��t�]�W(�J�{j��>����4�FX/h9V�oH�7yd���(������$%�P�U?m�O��g�Y���Q�79g���P��}G$�=<����H����ڄA�۞d�~G0 ���=�OQ��%A�z�*�_��(ػ��� �v�R��K�G��C�����V�{FN�����VN�Ӕ��������E����ȃ�5k(�Cw��A����S>MIRh�� �V�ڱ2m0D�X��ڒ�aX����'U�|��.�զνlP�M�C�FHo��m嗔�c0�2<�"����uh���>G�Y�ֵ��=��$h����ۏ1Z��� �����f��e�q9c����H��y%9]��N�Wփ;~���!2L��e�?*9���R�7n��@��L8 v�
N�f�@q�2�Lw%�H��`����a�YE��zn����p��ؐ#1��[��?�Z3%O�����yz�R���k�郚�0@g���L7�x�Ps���(��_�H�½�E�͸�.���%s_�y ��{{����P��C*=�7j�� ���y�׉)Ŕ6a=Z��^<����ZT��ޖ{��-�f	3J9��b2�y� �y���kn����1I�(�>�?	IFx?�DSW�B�����Twָ�r~��.v86� a�e�`0�`��]�b~����.�x�mDv~g��KVt8�Tϓ��۟��+c����W=�{SU+s3��!1���Bs�l<����DM n*��l�Hn�U�5�±�����*2�O����F@��[�n�?쨊v���X	,�/�
C����*��ߊ���fD{��/��Ho�\�ʻ|v��q�r����T�϶�r��/�ן�.kȓxTu�����l���6b�s+�K�9�4I%�l@��Ƈ
`ðmL����Q�uM��3΂v���2��hy핏���K��/],��h���A�qV���/�V��������P��prK��uUpǽ�hUe��aR;^|�T}�n�nF���2o���J�� ��/W��gu��x(��ض?n�@SD�Kc�E�)� ,?�OG�A[�U��19�V�ა?3��5�k��s�I��,x����W��u᨞���x�A�<�T��[��)��G��>b�`	$���ysH���@A�ե�RJQ���2_�p�
�f�.?'�ϡc�_!��p��I ;��Nnm��o����V���io���(}a�|%����t�ް2��ʆեX=A�Xİ}�o�����%��]�>§}�Kz���[E5��D1���(���u��vN��d���(������└J��3��s�Qbs�R%���;�ƛ(ap�r�����~��I@ќ�9͔��g��pK�[�`QkKS�l[JV�g�2�{M���Nw2�C��{���mƻ��J�?ϵ�+AwR8^g�,�N�L�����p���9\��9��90>A�]y�*�)�O$�4��K;��e�	��á�ny}��R�!���nk&�7�h+��D�H����i���c��
�������5F����y$ �`8�?�|��T�/ټ]�T�+����sֲl��a2
2.ӗ��!�ʋ�xFe��]�u�zF����5ܙ^�Ŕ���j3xaNW�~w���}�3X?��n�W� g��Jx'\���5��� ~Y��˻���#����DI%��C@�ih������T[�56��f%m�Ņ6X�r�3�A��wC
��#��غ�����"u�)����Gզ���u�e-Xz�2z��PZ��d�iQ��H��@4�n��3���d�(�W���-��ݪg��?�Cښ��ZGș�~j�+�����8O�`�G��]�ϱ�#X6������
�)��'T��u��gD����:i�oG'�PL+s��P��f������k`����=�X0u�;6��,2��4:�D���� q�I���(�X�~y{��U`4�P�����8s�O�V����=�G�1�4�m��h'6�L�;�l��}Q�9
��.;�����	�4��(9�>��{Ꚇt�G�y�p�.�R�Z�,�Z���V��XUvdG?�m�pNı����=����4?L5o�3A�.�Q�z�<��ASe��fE%��͝�H�����J�	����}K*��aXÂ|}Q�����Y�#V�yjhxʟ��9W�ZigyJąiy'������qXr�����;�Jn��K����n1��9vy~t���d�<�R(�ǝ�+��q�jɨ��7��Nl�"\�ȉ���k&�0�],3�u`��������gw��irx��_�������z�g2�t�����8�ߏ֑���U�PK�4@�Ƞ�ܦ�P�+,�C���ªru��j�(�d�� %��V)����o�2��
�hQ�0ko��s����Eܾ%i�s	s����H��'g? ����2k�t�b07���~̏8&E�������hc\i7���B�d߻��e;�!�a�ÅV�=*/
̈-�8��e��5˻���zB��pk��y֧���ퟥ���?��/@�q<�P�1�k%/��$op#p��
�ٲKo�ov3F-�m���%�}�:���1*cN{�ue���,�X��("'���LM�%z�������*i�7�G�E2�%�Y&�Il��5��8])�#!���
�dyL"R� v@*�<�FUvy�g�_��Z�	����a�o<�u�l�Űދ� �­ t���;᰷=�9@3�$�Dlz�\P�?��q�:Wэ��O����!���i����ex�i�n�	_�~�q������gnG��B ;5�N�-��B���w%����������3J��KG�X�5Dc47�&��Rb�E���1k�P8���C0��P���mف�x�"�(�� �x�8�d�Zys>$EݸG���ݳv�Ǵ�6����GBO��za�x�E�~�	o�hĊX�>I�'H��@���C�Bn~$���"�ѝ�[ޤ�J����r�F:�[=]�.\��&E�$��7��Wt2)�8^���0k�g"x�P7�1��1.!��H&l�P��-��|���l	���R�&s�1���xjR|������½��F{�v!a���f85��({,o�)I̠d�B�_��;J�g̔����X�向t?����Xp�<h�k?dsas+�cE���VŞ[�\z��7.]��C����ڷ��};�i��w7=X��I 3�j��I-m��Ù7�e��e����D�%A3����
���aq��s�"���ZcTKT�D�[t-Τ�?���8$k����: N�tx#������]��6��Oi�[q����fM����`�9�ÈQg	y?�	.(�@Oԉ��Y(�:�*���ǘ�|��P�P�60!�� ?�#����-O��x����+e�j�'�%m�E��߿<\��&e� �?���n������ߠ�jE�A8�Lj���2���+բ��Yw��
�@�.O#!��V�����.�L. �	�b����Zb�!.#λ���7>�#q�r�\�8�Q��
]�;�����W$'gq:���}�5
rR0����u��':���D��d���tV]�Y�;:b%_wM�R�}�>d�<:~n]�j�I���9�ְ�-7d�������*T�c���"&~������v��� ܻ��T�O�ʠ]q4%���R0�nL���weT_�PPy����X�I9Ls�^^s�dpe����lNs��`�֏�������k1~���R/Tk�L�U^��'���k$��Tj'	�=��T�[���|7�1�bS�s_����x|�f�d�mE�,�w�� #��2ݤ:48X
��"��0�C!(�#��|&֟L;�P�=�uh`;�p�dO�'���[�&�%ĝ�P}�n�1H�ߛ���p�����V�dk8Y�6�ŉ��&�ilrH5��5��ѾR��,M��3��F�z�lm0fJ �������9�e)c搋gdv�KFOnµs�J�`"@l�9W-�,c��g����x�`�ԋ.�䖀 �;ې޶�R�Ր�:ӄۂ�!�ZH_8W�>�(?uB��UE��i^M�O%�1�d/E6 ;�+(�=<6��^C�}ϭ��Oh��E)�F.�g>�t��J�*� H��0���[$���9���p��f�}��C{#�Ň,��?q�*���?�x�䍵
�E�|K��S� �V�f���|��툉e}�a�����R�&c��f��w�W�!v}L��
��p1-�+FyE��Nu�z�`�Ϸ�"�a�7�ﰛ��,�;�`�rx����Nw�Q ��y�����?���bEӴ¦(�Ku��������o�����o��TL�ٷV�������ikUs�|�W�����/��b<a%cqX�9-h^:���,�{gGuދS�!�y�Me��ֆ���,b_��'����xԹ�Wv�G���]�YA�,b��� >�d�"�Xa,��M]�����3җX�`����ַ�<�Hh��F	��P�F���	�RR�,��CS7wԁ뭩���
�[%��@�{�S��.l~lJ����>���0�q�a-2)CN���\��B���W=y�h��j����׉���'�(�vώ�7�:d=��5��N Ol���y����L�0^Y�
nH��h`���@�$β�b�T �J�$i�ݺ�J�*⪖�7�0�R �u-$o�H��;�7̾T��}�P]#�W��k�ͭ�p
������q�דi-7��}��UT���7E;"����kV���"���g�N�.��a��un����p�>Y��a^���!eN�}?�ؑ<)q$p{�� +�L򍓧�ȷH�g�=w]N۰���3 UɄ1��W7��5�^/����� 8��X�,�r�d���;����NdiQ�Ћ�1�u�w��\������9Ko�pV��X�q�|x}QN]�Q�+K��<zNW�f���5��^���l������&T^��T-b���݈[�y/s��5m[���l��;����|BZ�o�/�O/��B1jwEJm	��nz滀� �W$�ё�*���Kގj��v鱒�zvs�A/�׷*��>B�#✨qK�|cw��rse�,�۾�P&N���IE����slU姰��q� 6e3Ůa(��h{���U�p�?��$���e��g���U�3&��� ǥX�U��e;�GLܧXɐ],�v�{�8�y�^�;�����b����/s��Y�w�Bx�til�^ҋ�wd�8p�g<�xqJ	J�\z�F�m�y���W�!)���h�[3qQ�f9���t}���?D���$�Q�x	P����D��ȭN��>}#|����� ѝ^'��87�O��7_0d12@Q��}F/�C{�,�20�R�g�E�Gn��t�Uj�<t���o��i���H_d��Y�~�1@��n28��G�0_�h�`�G��)Y��.��F�ր��s洆K�t��]VWw.�H��(n�	�,��A�Uh�fwE����'���g��<���!�O����z�c09V�����潴��G�3��8��0�0��9K�	  �*q �4�q�tL��Q>J?'a^�I[(3�)�b�w�^'l�ۜbc�4�p,
��𝃞���VG>v�2�Ѿ��Jshk`���e�e]^���x+�_��$4>]3z�H9�F4��U瓮nc�_�5���nP9��"`�P�B��U�v9�n���h2��fN����c�G�m��������r%h�	�1�r�՛p+�a�%�3�y�9[PU���ǽ��;���?(B
�5i���x�WD��͘�O�gm�L���s�=�Y!�^�'�]ކ��Z�+�"������G��\$h�E�-����p�����(��I%�s�F�줚d�~���p����U�|�U"�f���)��NW\�;��x�B�l	]) "s}���3N7�+GhcXK��3��d�1@˼�P6j�&�0հb���G�Z��l[6[y\莤�<ｘ`fQmW;�����b�_��H��x�U����M��A��e�E��)����K	2���8LM9���13,�"�g�7A䞉Z�:�=b�Q�u�N�C~��"ʻP���h	C�A�ul�
�������GɆn˜CV�M���<`X�O���#u\����MH�!86 AUc��u����Cg�`��(�! �RHA�D�x:(18����S�d�	���:$*�V�A�a5�/�.�#:�(�su�9���!֕���X�> Jc��°${5��o���F��`Riz4���l���g][KK]�^d�]���s�x�2'��@�g�Y���.��)�^g��=%|������N9"�?�s�(���]%�h��=L{AI�s�\�L5���\P��T;Ny`��HX�/�o#|��G8����y<�@���6:�H�v�������7J��nw�[M��F���j�D�`�=���4j�.�eK�{�z�;N��h'қLY��^�� *Pruí<P���H��H��a�V�IK>��D����S���L�� QVb��ޡ\����5�Q"��}2��d�d��I=9K�855�W�2Uq~�&k�B8b��y��z�_��̂<�ݚ2�e.��i�5d�ox���m�>:���y��vt������d�%n����S���,r��ذO��ő`���"�73�4�%�)��3��s"�+�����o��m*J���Y/
���z� /��*sM��(޻�{���q1��5#�]�����>�N`�����˕��N]`ӯ2�f	rPMz*,��_:?MՇS��S�T��[.^eF���b��:E��a����R�Y���Z������
6X3+��D�e/j�R����0o�8'���f��o겂1'X�T/N���d�#k����EO���&�����'W�� �:6���G_������C����*�L*/vD����ځC6���1Y�Iq�ߌ�~����0��3��g���m��<���Ԭ�ł;�M>s83ܬ��}�b�̓����F��,��s��UD�/�ｰ VEs��.lt��'z��F´%HN%$j:w��ၢ{�Χ��G��Q����A�m�zw#zהȑ���|DId�z=˓���y��P��G(NV-���(LP=�N�.�9������i�s����/?�-��W��CktS]f�U��9|\Y�e���H���ITAR����]*�R��U)t�yM�	�[%K�W�_�����o�{?����^΋�*9��4N�W"5����h�-{	n���bվ
o3pa�ZZw�z�-����s�������r_��=AU瀵���2�X�eo�����k�tǵ��*��y�3}K;x�#I~�"ƖM���{Zn;q~��'�������Y8�Û���ȫ������a;e�>^���4��Ů���t�ˣ*�_B^�ߡq����n��.�����q�+60w83����AaѬ�5σke2;탏�^��_AHa���qPuk�A�(�x�N� �hX��]ܺ�5��3�B5ʽ]�ί�le6�18Ø���r�@�蟉�ڤQ���g$�����]��}o��<�K�(��i�en ����E����{�r�v�U[�����,0j�jD�6��N��6M�R�s�OY5EOL5��ɕja��Y� �| �ݤ�>��7�С�˩�R��=��Dݓ�OZ�8v�j�S�7�������#����]�[�Y�a�3i"�[������ᦑ���25`Sٿ��/k�픻�H���� ���S��pw�~�	W+K�����^�gi�%�̕cklp�^����W*�R��g��y���j	P��C�&|	�6�,�?B*��vb�-���r��,��8yW>�c�Xx��T-�C<�[�c�É182���\ajF���#p��T@n �>�`�U�,~��+xV���y"�sr���Q��ҹ�t���4/8�ϛ��%�䁈�"���2��vlp:Q]1.�p�>�K>��dƀ��;�܅�����@�~X�� �������.=�$/�
�fN���=*Q�n��L��R*��%����ʦ�����G��J4���T����*�)��ZI�CF�yu�a�cSt�^��S�A��_�B�\f�Z^��#i�-Z}*�66��GpK��JD��"O��b8ț�ZGĞ�!��T���#�%��SlEn��P+���e�9؃�����$��^}ѹ�P���-�j	y��\1,m_w3�?w�Ӳ��O�[��*����e"��Z�M�}�n�1�K��@�@Q�d'�jj�\�o��
�P �ˌ�O���u����}v�?g��%��LgCC�*5pаƕ�-n���L�L�[wX�r�>����8_�E�;��
8k�Qz�q�8����);Aį�v��F�~�̈́W󸁟:��ו� 	Q���HR��xٔ1ۮ"(��^�箷UNjj���Kq�$�D�@ӵX�#w:�,��&�z��L7A$���1���9���4����ˣl�*���[]p�}�q�P+s)��~hCSRI���%W�%H�vN [�4.<����g/r%P�9_����2��Q��,ɡ�ptfo8T�1G��v�Q���de�F��)�]��RV�8y�� �,��+�%oO*cc�����wM�E�R�2��R7i9�ip�N�t'ާ�ojX1�*�]�5�Mن�VQ�>_b�@��T�,V��(�s��1~��j�6˲WQe$A�,��0�)���>@$�>+�Bq��#�@i�?�<�>������z�L'�����ʽ��;�01��
㞟v;C�X��8%v�iG`�����j�A!�#ޒ'�{o�mԂ�R�A_����p�,ZbM�Yd��^i:��n������6��G칹�8�ʌ���Ͻ����H
<n�@��M�O�>UK=x	��A+��P�R<Ӥh%Zr�|3:���,
�kh�tsg�X�*_��'�5�D��>�פ5
@5���O�ȥIu���ȭ'x�O��S��{��`��pËH�$b��
+x:�S�dasޘ�*��b��T�}S"^�̛��h�j����
�\���M�o��
RK�͛���o���M81�Ԋ��$�6�����~"!��4�1�R�͚��I�I�]|V���eZ¹P� ?�v}�@5b"�MS^��9��/Ӻ�Sh���B����Y�*
e��~����� �DUn3Gn'�7��N�uG�×���Z�ɽ#��y�j0
��ۗ�eG�S��^���c��WY	r�O��"p\!�pq��Ȫ+�;�n��W�q0&�O��|`���`��;�j��W2Д)-�l�����.N�?�ú3Dqt�>����Nr6(g�=�d����H�߻��@�A�z_Ģe���#���Ch|j�f,�51��L)>�಑��x�L����]*��͙ y������/A�Q��qO�fH��\�a�3`K2ϻ+�v#��V����c@)����s3��Pɉ��C8�G-l���q�\s���7A�â���f�uha�e�h1�DysɅ&�㓭�:�#�'~N,�p�R05~k?]���meLf�zi�t�)���s�SQ��t_���M���"��5��~Q�Zg��!�qOZ��S#[����#��8���y�g\_�������Z����و(vx"���릀�%�eT��I;T�J�k\��"�]e23��6�^ķ=���f��:�}�[�������s�*`(�(���oΎ�l�mQ�`|S(�o�F?�h.$�v'�O	oF#[�R�l��$Iȝ�G8(?��i��nMAek���5�Š����Bz^o�M.R�����)Ó� �����r�G�Q��� 2��#�X.B��WXe[���δ���S\�Ba}*���
�H{8�:�������C/-���BRB����+hF��~O�4
+�Ɣ=@��8����g�!J��J��;�}�'��Y�q��l�8S}�Z����sp�N��y�� �<V/��H�٥�<3a`�*`��S��/���	����q���
9�Vh3�1���x?�-�!����<��� 7L��V?��8M� �|]�����kI�8�.�҈{�cI�si���	��޿�?@��+�_N�!C�56r��׵@�d#�Z��ᨭN����!�q_�{�Է��4�p��5�Vy��	���o߯�xI�}��u��x4Ue��Z� 4��O�'������l�/�G�4:c�<� �{����<��%j'�K�p�q��8�0�2�fŏ���"k�R@���M�U����>��IM�}>'�Ds���o���m�[Z�f�!�2ܠlY��M��`MC+���%�'�VP?,���!F}sD����:ô+�`������@�L�M��
�gG.ǵ\��\v^v�h,l�|���1�^ҋ�dKf����z�C��:���fJ���It"o�����R[�%��W2qF����t�&О`�!PFwb��`�nT���R*�(�)�����MZʟ��#����]�y/�QR[�8傪\������@l�2�xm�M��a~�ߘ��U=���_��)��vY��#(�b ,�8r�6�r3���w+x�
g}��Df�܋�w���uL����Z�dӇO�뉴�p)MA, ��l����=��}�d}� ۺ�����T0�]�6��b��4�Y!'1�p�����Y
�m'6PG>�٣�W@:���N�7B�BT����bje]�������8l1[y���$�H�Z-�Ic���zgnxXӒy�tB��"��Vsȇ���/���L&]1�� @q�<��7�������)�*���Ai���O"�gR;�q��?�<�2l0�71��T�_������؊�����p����'z9�6����L������/����[}��e[�9=��vz�B;��#��,�jc7������L�{Ӝ����.���ٟӥ�LP�1�f2���S�Mw굆�~ܢ���z�'�_Sު?����Oq�v��s�{w\%�k)�k�Ǖ%����Lm.��J�P�u0;CU���ǘS�n�b�o���A�������cC�z�4���ǋtD�ИG�ښ��J� ��W��BB�&î�~V�e�.(�ԦBJY��C�,-�o�N]������k ��2[�n�]8]^H�oU�|�E}}D�����8F~�E��>`A�&�U[�P�x?ɮ3H���O�·��mr*��F���Ĉjy��綂���p� �����Xy-b߁)Ԕ�E�8�M������A��X�3/	Э^O�nf3�
9B%kTM���o|G�D��p�'ls��j-��B����
�s�����@�vꤿ��߂�{K��	j*��u��)�����: ><���j�Ҁ1
������b�pFQn��(�YW�0�Y�������L%�+�d��>S�+\-ʦ�:����ⓐu>R��3�t�jy���¨w5[�25+��h�X�*aӕB��� �_�*諲����*_?�09����To�c�!������#����,ypmT<΅�>$X�T�L(�S�ԧϓ���Ϛ��\�0W��MUO���JLQ3�Ӵ#0J�Յ�r������
�v���S��&���n'U$�4����Sb��
�d�	΋�ݾ�p��K�5�^�Q�2j�i�h�/��Xq��2N��4,+4�_g��_3;��b%�g+�S/��\y���oG;�ܬ%S5o�Q:� (/n慠��+!n���$k��ʥ(��QňȎ�>�%�+�q�\y�)4�v;�1�*Yv��7q05�yH̓��@�=�1�����ZR=�t�#�G=5�&,ya���e���E�7άx<d2Z+c!p¯M�1����l�Kf)��6a�܈����,6�y8|G��5�h'���jĨY����[Y� ��$�څ0�~�ݥ-Q-g7�`�:�nJ/j�h�FZ�Ջc(���Pa:e4Ý���E�7M8��e�`R���i�0� �5�#U��k�!%�<�� �o���e�LM�<͹����g�����+��$�8$�� e�Af����z%A�2�da𺺳��@<���^�DB�ܿ�����U�P�r��;A��-%ב���pK�$��'HR����P��'~FDn�꫘��e�Ű�[���owOL��Tqr�V��Q����k&G��W��5���9�o`B_����`��(ݸ��!��F����OH�C����4�г\��*����ZW�����y�Qc�&+�<ܰR���A#�ҔFA�q+?m$s*�®y��
R�2�Eܴ%x�ؾ����q+���
ۄ�c*H���g9�=��R�#�V^�e�h�/�	X�V�l׃��U�Y�9�s�����{����:5��v�d!y�R�	�l���T%�5+4����\*}ƭA�-MXFN��lt,�jBP4���U���y�r@�*4�ڤ�Đ,����zt��i"��-C�W��g	��b��Wl����Wb�߉M��$�#�+j{V��z��n�C¯�5��F-�\�6ҧϾ	�f�K���k�?�7p���e�xD"��mE�*/�	���Z ,CX��'z����p�i��@�|r�oFeQ�j�r���˿�������o�;�\��%2..�~	ojO�bɞj�;j^Z���U^Mם�%Sv?|�CBH1��3�.���O�׌S\D!�!ҳ^ɞ�@�s"��.���x��5�j�����=0:/gjv&q-��6k���D�>�s�K�'�jd��HBx�H�uQ�<�w�N��Y�yG�ZW.�m|Y�4Y��7�L�dR�P���ƿ1F���%:�f%��ml/�z��V\���H�{Z�;�iH�~��3���z��wP�̓J�0ڝ�}�-k����q

Ntd�lK�;\��<߆cI��:�>o��VZ��>���y�5nKR]B}ʬ��>D+��)�/�y=K&��f4����6�t�����ɭ�R�[懕�m�A>��I	�ݜ�'<�&e�=l�|�ï��u(���jM�(����k�Ԕ(�zm�ޥ;�i:03 ��r�z$HjXq���������O4n�Sf̽��l��u�}m;D�R���\�����ǮX��e�H��/�e�Wp�,r({���F��y49�;��&A֭3�Hu������Mͯw�w*�"�uC`T�6/����Z��pT�=O���̗�a��$ǚ�`��Rk�d�>eΣ�D�K�,�y�*xH����'��̜�5����!��-_Mh2�G�s}i�V.�ˀ�l�0�\_��5'�a^�N3[���_&��1>=�#(���W��Ɩ�$��p(Z�q9B���f[��Zŀ=E|��TX9ʘ��F<71����=�ox�14�At?�N�YS�J�
��-�G[8.�E��G�?����5��w�8#g&h��y��+CdPձ����_��O]��q_��=��R��v��*��� ��B�Ze�����-��y~x���� ��X^���P�¼	�Ӄ�����s�����ݘ�M��� [��*ڳF�0%������0��ʩ!�xꗔ��u@���Ч�ΔZ.Ë����1��nD����f�ޔ>�^�Nܒ�ҽφ���e���l���I�	��������y�����py��i}|�x9'�ک�]�n:�Z��͍�� W����/v�'0��{_z�f��C`?k�\�bȹ�u�e�����q�k�^5݅�5�N��n��2hV��{�S�/���c�6���$�5}ztɗ<i �
��@T��I��d4��A>����@�y���jڸ-������zM�&�}�4Z��������S��K��E.^�!`���8���K��;���!��R������/Y �o��O�����~��G��#yo꼦s�� �C�ROA�}].}P^�M±��7/��Ʌ�좀�w
XhQe{�M�@�]Y�����[W�>�=}zƯ�ʆU���נ�j��bI��هA�N0V� >�S��D��_���=v�v@7ݰ�@�	�(z��E������+3���Hp:J���tU�O/�f�4b0�y����I9�t��M��{=��u��d�4��I4�ft�8����'1�������:L,!j0)눷�D�Xs�ٲ͎J|�L�S�f��Y�7�|W�.�/E�I�Uu�no�h��>'{���Ԙ2�qKP�5�c����uD@4�!�X�����	�2���/#}?�Y�-�=�g=~ZOׄ�uM���;��!�|��v��6��҈����9�5Gɻ݅!�%����d�.�|��H���2j��M��&*�V�����u�}u(��1
 �Ц�㙳������D�Tm�&m�y�^M�A�W�ѐ��@Ӯ��]b0�g�g�3����6�܀�p���9��T�� je��O�������::�����������(w�S ��Zux���~�e$�W�;RY��$��g;���3�z}�~��������e�j�ٷO�xt8����K~���%t`���i��4cM�L�#%[�!㇀˼���=p�X���F`>&�Ά�������@Y�'m�03��qn��#{s�˲���&�H#1}���n0�D(ɣW�xDwv��E	@�1���ǖ	��k�FxM�X,?�c�F�''L�c����:���@�_s �L)m�H.��W<Y���P��w���%X@.��|���Z�@*�����쎘,�,t6�����a;�N14�I���#ʃ���v=��vF#a�s��;U���9�K�� ��@OrQ�L����1��A�s�n��1}
�ڶXJ]�� ��i�
y�1��v_�\� �}����[��2qk[� V�8���Jɹ�ʑ����M?������lsfT][���zv*�4� �:�]�l�j'"�mEc6��
��}�ƶ�s�Ĭ�[1w��>���z>4IsJG �POb}����岠j|�������UT�_�,��k�\k�r���o�/&[־��Rˆf�a�]��cc���s��D����c{�Sb�N���d�S�6Ÿ\R��r[me�;8��yWe��}԰z��Qר~��?����q\���[����9�Vћ_8٥�Ao��� Ɖߝ�]�{���`��Mc�����#������R����)?������#J�)��XQ�lQDL�>����z�r����C%n���D��3��{V�3]ȉ#����K�t�
i�4�K���Zu���?�ʰ3Y9+|;o�{Mm��0F�� 4F-wK�1� n}�A�e�
h�*ST�b7A!&����O�I��P��X����l��ϼ�Ĳ.�ۂ�´���s�ĳ�g%��z:O����n�"��#l���'����T�kR�A��@R3��n�#e�WT�����N&�_|�gخ�Y��I��;�l���qT$ĩ����H��L���T�qv���W�iP�O6ov�zu0��9����UJ�o;ؽ˕��|�B��b8�z� >�lbp��Nr��#,�:#�1\E������5?Y1q�#!#�k�-ڧtC��Q�hp�8.�r�=7������V�_wa��:��en	w֬ä�[(�:���0��Z���|�����+`�D�S��QZ:��Vh>�E��j�b�� ]�} k�Z;A'dJҘq�=H���������&��-��e��m�*9�bO�b��PP�.����A�!�&dp��_ �yTp���1G�ܰ�ؾb��GyK"Tzu�1�UfR����R����p��T7]�[�AB�[�k΅$:T�1���}Q�^�hrH��kx������gk�gW�F3�U!KF������*�l.#Yk�~	�t�p�ʮQ�N�س�rC�4~��=XC�Lv�_l����W�HB�4��x���;�*7v3������%n-97d�h�T�Z�?|���mZr���ڧ���J4rb�����$g�F���trf�Pq��hY�|�:I��21�a�u�`�#�d^,T�(�jϥ�q�n��\�f���D��*x�dzT6��6s݅X@u1*���J̊�}�b�߾>�2R����?�I��)���+�:���a\\����Lٯ������RY�������&��%��t�4�(�Q�N��5�6���%���ˑ���B�]��y�ےo��Q��좋b���(}W?�vP�8�)j߬��.ì����S����ed2w��e�X;�t�i҄�=�H)瘽����|�f���|�� ƅ��*��h�
h�G�|���x�؟���u�:)�Ǐ!�s��z��8A�T�(��=�������3&]��7��&�0,�RD����n�(õ{G�J�`�{�VR�Qp�yZ.�?�1I�����9�
����h�]�AN��v�e?z�u���G���F��x�f�c}� ���7���O�W�Ny�(9��k�yD�Б9g �r�PhG�O�O�gxC`W�G�]�;�*3Ⱦd�#�wD(�N_��Swk�}ڎ��3$����tӳ1m��T����!׽e���U��,�����l�d�u6֋�ζ�H�úq�Z��N�i:���@u�#U$�!�	�V�GX�#0h�L Ȍe���7�~�+,A�J�#@�r���Y4�r3n1]WK�5��,h�{�8�)�>��	!$D�_r(�b��[OxkP[g��×��s5#B�J����v�W�%'qܽ���m|l,��V�|�
J!���h	���Y+^�ጿ�Q�x��6W-ȓ�><�q)K�F���`�۠ƽ.�av�U�"8�.]8$~l��6NL݅8�~臔��[��E5^�S5�>$h��%���f� U��A(G[D �]T�r�7o����}Z�GN^/Xԟ���ĩ]PWEb�" :�Fȸ5t��OB)
(tR7�,�Là	&�l�Y���-��C�3�i�j M�ř7�g.�a9�5G0,H�wZ��������G[(]/�M팇��G�q�j}�ރ�~3<�(.�	щ�Е5���$����K?��X�a]|o�YS��$>o�}a��D�l�;��}do�S����j}ݸ��;�:u���ӎT�'��4~��\�i�!lX�C_{#Og���c7���%��%���"�i�Fy j��?O�W�Xԏ�h>�_�O�}M�1}�l)��g�"�dr`m���5�"z���/�uث�wL�P���
�"��:�O^g���r��N$�sE����y��G�~�7��zo$3x*ڭ�LJ�0��eu�9MY7�پ��.Lh�>����1����i�	�<E���XRnm�&��eg�<:upq[ ZI��c�%�����+�ƜY�?�U�I��������oq��u��9g}�|Fj-
'.F�[�06mD�ã��ԛ
v���s����\���;�c}�B� �v1�>f2
߆KE3͌:G�t��{3�:� $��2��?���`V�4�ˉ>�/@��R)maS��p�B"�M�␶#@�/t��*z�=w��[��'I��M�]��ӀX��H��>��n �Q�Ԡ�N7��E�g�,#	� )���Š�ՠt�N�Ӧ���_4�Qю$3t+s8$���������Ͳ�`Y:� �C�K$� P���BD�)�,P��^��S9]ϵ0���X>gI�I��t^	�MM�:�|fR�YԈ?x�&UKC�e;���i\�䖖�E�`䭍D���lp~�"PEF��������aWC����*�_�T��̻�H��2 u��c�dn�)/:��>�X7�Oa�û�xeu�T�Ii�j��xV��ó��2j;�9�0���Y`��� �GU�P^�b)O1j0vH�@Bb_�=]���բ}�q#j�L�|9�<M����.-N�.ބG�����Ռ�k7wD�S����\�Q�ȇ��u�Q������L�`Sb�3Z�G��GN&a>^S�s�KLA��X_a���3���	��Jc��!���z904����X��L�Nqn��� gB�0ѭ;9��k|B^{���,4Wb�A��MӮ�%�'�m��T� RJ�6qOF��ϟ����G���nyߥy@[
�f�^����R�1�I�fk�Pq�,��wZ�+��e��h!b��,���л�Ţ�\K���+�')�^�$T 9֑���^@���i��\ ���P��l�f�o�cW(8��(#<�&��q����= H�t��_��}�t�'EJ\ڈ�R��\�k������n�kx���$`�y�j*�*y�Z9�ے�s�S�hFl\�Q�9o2��i�<n�6��)�ں[,��Qζ� HN���Y�J��m�n���Y��&F)��+�[k�{r���z���M���(�C���:�[�[�j�����+����`���i��L99,߱�,�W��]s�&��H3���U��VO�+N9uckUG���R����C�eU`���}-��ݽܥI$�W9f�E?�����5ŝ6���U��x�(�ώ�>�%M�f{>�$��4m���
C3�Vg���Mƙ�eݓ��c!��f]O��[ۀrN]E�̛-����PˈՈS��.3��~��!��٠WE���hi�  ʬ�� ������1%���n��4Av����L�ZR����(���H15Fe ��i�@�W��L�i�l&��������l ��_�O5�PQ�$F-��~�B�h�z~݃�FgȰ�A��_@C����6z9�gA��v��&J���顰�
�NAe.��Z+�Kz;��c����� &���M�ڞb82�M�-�$�e9�$�3��I�7��:GȰ �\r=�Z��:i �e4JԥX�F�w����s=�J*e�΅�gG2��[�����+�{'�r�1V���������.��y���}s��2g5�%i�:n,[l���Ӳ�"dͯ��Kщ�"c߄?����&�Đ @ڵ8��Jd��*�5~!���
ߡ#3!��;����S��s��#A���%�oL�1� p����\�D֧OT5Xg�Yɫ����&�+�ê�x�Ұ'���KW�nX���/���ҏp�������u:gQ���w���f�����+&*�j4L�6d��y��{���������t>�9����I��8����'�p�0�~a��Ks[�gtJ���``��t��͙e6�:i�KF�a$�v@&�������\��Y�^۠q������x�JLD����[;Sx.�plHN���]�Ҭ�u7gY��o���۠�*(�uS��Q�*�m���� ��?Y�`\�	�e_,Y���j��D��+�I��V��ʒ"�c�ӣu3��%/O�F�7��]�@���h��oD��W7q������KW�� �ZX:� 0j6�}�m��L����3�ɿ�uy.f���g�'[L��2܍�;P���b��2,-}��R��1E�,�2>On��H��5֛��偁^[�nX�1���sTC}� $�Dj@q��I,Br�h�']�Ϗċ��|���g��U;uн!`�o6�hW�Y.�'����{��Pé��>���0j�禩3D�;b�O��Y�3��~��F4���s�r�(�*�_�����]:���j+��7�=U��؇S�)�_���-�(�^T3�x̬�h�O�y���X���7���wPX��������SO
�+)Va��T�U��d U�Y��n)s

^,�Z�DJ�`��L~sU�l`��"2�<�`c��9HG&�-���~T��<��Y�k|�}JZ�?_�^���r��!\ߏ���8�����������_��.�I�F0�������W���`)xחQ2e��MP��������cpec���;�rg�¦N�Vr�I�{�J�^�` )&�����W�UlF%K��x���VV����k| �V�<���#�Quto� P#���1�,���8{��8>>WH���;��U�	�,_s7CW8_����MT9&{�(�@w1#�i!��Is���v�LTy�)��@�lͩҒaԎ��eV�3�M���q�8~]������ݻ �+c�^���Y?���m�P���b�>�7��t�޸�ڀ��)��l,qpb�+��0͞�v��́��]Tf�.�o�y�M���A�qEJ�n��s��An�u��������`����0��@�{�adnݷ��,l)&���<�$�k��Y�m�P_���IrXQ� Esn���(���'@Q��CӋ)�d��K��F RJY?%�ζ�dX�V	f*�@M8?�H2�S�%��5WM��lT:!��l�Y����|'
!� ��zu�G`�	5����@�ZI����^�����b�,'�������>O���Xlə�\�_Hr�q�۴7�,�(��S	0A�1�N-E9h�w�V,�5�J(Z'��9;���n���[�6퓚�uO5�5�CGA��odC��k�m�_<�:��~Ľ����u��t�WF��L�Ğ`V�>��[*�!N���T��}��N`�d�G$|Bſp+�V���/���&��WB*C%wҫH_��}7��0�[4`Ȇ�{��s��{�ːO�!�A��>�wPV��e���&{����%����C�x$�Ď	~L���a��r�� ���*s9�j�a�Qj�)� R=t�ut���C*��$El�}�0���@��-�2�7r��ȃ��c�~ߩ=4��EUP1�چ��C8N	О��A��K��)N�M<� {i�C����t��������z�.�|��Z��εE��V���}�.��������y]9�:�ӑe?=�)nOB�kq^~��!�{��`�$��U~��9-�d��Ә�Ղ�;0]K��azcs���j�1qZ&D��whbC�����}*(��L�nJ$5.�%b���l�~%i�5�W���8Dj9;��̩�3~�s�����*I�����>5-�3֓My��K�Y��z1L ��:�R	-���!)Թ��l��,�R�hݾ�q��Ni�J�a$�	�LM�gS/S
vd2Z��t�����g�3��Z�$ 샮Q.|F~��&�vЁ��5�Q����3u�mD��հn��[�?a����.�㦃�A�q�$�b+P5T��4�.J_��K��q�g��Tnf�E���7���D�����{J��?����%s��]Es���Ѩ9b���aP�۰�"���\�n�3�Ӻ\�ӑ�c���a7�eN\�vB&yh`[,B%�3��{�z�.��tU��͐�N� �l�c���8���
��Z��!����ʧ��*��d�Z</�}�M��~h��~D}T��m�Z��	֛el�;9D|��>�T�^1-� 0�l�K(`_ߴ��ֳ��|j`U��1f���vUB��0���&vڨ	'b�$�V���,���f��M�}�o�0-"�$]4�La���G��S)F�&����A�^I��`X�c�N�X��m��ȃ
-�g9���O�i5�+�ĄaF��E���J9���3�E�����/-��7Ĭ�xat(N�lZĔ�_��h?�6L����)Z|��%0�m`q&ٮX)�}`��W�4��5���^�����ˉ\ �ҧG9��\'�m9M%��ˣ�_ӟ��k��;�:mY�Z�`��ȹ6;��{T����"3b^o`L$����{4j9u.���'؇�dI��֙.AKr�h$�݁�Hu���)Ѵ4{�L��H^�ӓ��~G-�=��1>oS9�cZ��ɧ*<vp�}�ˡ����j|��A�j"+��6�����:��)H?�g��w�Q�Y�;;I��n�iz�%|�����&Y�:��Ay�ֻI�������;x��'�~�3�]�F�Ǿ��m&�gm&P��ͼ��OJ���֥����s�ڧ ����u![|4VM�R��M��H���J��{BD��|=��p`CW���S9��O��98���8��\X��Q��I��.	����-H5~B��/dv�B����	֩�\D-��e������X<]�Ǖ�/������_��9v�I6^PY��y��q&]�XqjKi���䈷�yz%��LS��q�" m���"T���kF�,@T����ELe��&���9ҋ�8���*a�A3d�l׎���e�T�o)GxU���6{r��y��\ap�Rx0H��аv����)����\c'|Tփa�R5��U��mr~�s�o�|A��ܑګhJ�D���������2L��yZ�/Y�&E�#D���4a3ƾˠ��ۘ̄Wb_�h�Ѥ���\��w�|�����]<�`w�- ��{^����=�+�`�a����_�x1�����2�s�´���M����Ʊ$�A!]�r��;Ʈ��@�	����d�ػ��O����ǴBˤZ�k깐�O0v�ҿ?	�\j�al�V�}c�+��l���F�=��狣퍕�a�qyN��l�L��1�=5)����d�tj>��ޣ��:�T�e���z�Z�t�[f�N5ڹ��K��'����;)��zK�ԛ4���u׭�d	�(���C�x��RP?^��CƸL����\�|�v�@��숟� ~IW8O��]��wO]
Ȟ��7��|�ׯ>��/��n�p���45'�ҥuΑ@E���O2ܘ���/&#AB�Y �rE�n� Х���5��e�p��A߾E b��SI�s��A#�Ѵ)�&ʊ��;�|�%��'���	��Ej^R�0��m]KD�{}o���z�L�}+�q?�H����yuZYlԅR	C���I�02�V�s�� �)��FE效�P�����7��0��r�]Ь���_�d��M�b����s��~��e��qphi��Ma5SE�/ݚ$~��U�(n��7�8V`��Ho䤩O�zO��jS��GD(㋍��X��_v������Qe�.��6#=����m���s^�U��W�\h?4Zi������j��&�ڳ4���(Ę�6X���tA�SC5�N	�ܽI��JY>l��`~��g��Cb�
�;<.���a��w�
F�G	�C���?���f&_�w�̵�i�I)uw��o���EWC��2�9"ĵ�}>^�)Nx>�����Tϛa��aI���j3�0zW(�L���$���p�*�����N�q��ɜTW�ٰ��y��N��6��=*c&B>Dj%i��HܢN*��|�E#�������̭����C�()�W��g����\L(�]2��9ᆐ1�ݣ�hK��8FA��B}��bL����$?2ԡ� .%�f��&���9HVw�[Q��S�&��Ҟ�Wx�:#gm�d���-���YaVt��ۄ��#Js���t��H,C�Ьx�mĠ�1!��0㏺� 4��Ѱ�Y!n8��C4� :�"�.�@!k�c�<*0�&�C��ݐ�W@Z-0���e��ȅ�K�?(�]�2kM��uB�	M��B���v�
�����Q%�*[V�T!GKJѻ�ު�^>3�r��a�Eq���1g7����h.�}9@@��]�[��I�J�V"Y% Ǽ�V7��z��f�;���j�&z"g��C�	��\�T���4�=+=�=��uD5ye�����j��Gڊ:��������tř�2|��z��k�G0�LwY��0%�II�ϰ�q *
QJ?��`ep�|���=gs�V�	0ܼ�K!C� ��5$�QS�� ����r5��{N�H$��DB��
�d	��4=o�h�5�՜v���H���I�M^1�OU��,@!�}� �����J��l�G�!'�xo`Cx �b�n8�owZ��@p!w����	�u���F=A�����~Y0�|���z'�rJ�%�A��¹��`$A�����v�)T�Cw[����4���2]_J}��[0���Y���`YM�y|���,�^d&a;˰���)j��1`������t<n���O��Q�q���mh��X��Z�4��=�<NTq$�:n�{�!���9����E�Ϯn�C��1��by����Y �
]��\H��2�Ul~�(�хSj>xx��U#,�C�{�c�X�,JW�y��I<�DھM�k�^I���(x�p�*�Ctg�fLe�1����a��_��>��.^������fD����f{��i�+^��h��ζ�n�s�p�~����+Ǒp/K���<H���m�+���/"� ��E+eME�{z[k�4!n��C�e	Y�#ɸ�l`A�-�����6pZGK�Y��۹��i7֛C虎QOM���1��j��P�e±��?�NP�� ���D�.�������w���W�D�-����"0W;X�d2�s�����t#@�2�}6<�K��Na�֭aX��l8����	J�ZFF7/V4�� \���=j��]%~�M�.��)�2:����K}����Ů�w��`!B����_��E%ņ�s����@1�"SY��sS5�u3�=u���M[�e��!�pR�@����)�;Yq�>ό�&[B_5�I !E�y�t�sڮ���}�n^�}`f�d��b.Bա!6sC�[�E�p���>tO�ǪT��?ֈg
�k��ճI�P��,���3�f�N�s'�x'��R�&���ɤ��+��6���G���kr�3����Sa�^Q��ѯ��>##D��Xk�Y6��vM����W�t|��&�beN��?���s[@6q�``<�S3y��c����.V�]�5ڀ�Ď|5Ԣc@�c�����y����΅��b��1���)1�p���	j�C���雐��#)`���n^�r8p��p�3钞j^�<���������$S)�Z��"3�ףx+���>�0��|3���~����C
T0�][��K������5�)q�d��� 9�m��D�4�;G���hS�sb�y��7Xj�x���ei�s�]��~�]1y�+
C���2|f+���Z�[�a�묠Y"W59�Q� �A>�� 0W*����̉����5�z���f)�Ո~¹�4�i�=B_!j����~ �x��EbF��ĉ�B�%�Rb��%.�b�S�p�֗���*+�@%(+Ng�dt����1���ޢZ�}�
����va1�p�%x_\��^K3ݝڛ2;��O�M?9��C��;����Au�����q�7�Z��W��І�c�xzN�Zd�] �Few�q�l'P%i���AX��)/��߻��r�;��_�P,�׫�5կ�3���������g�p6���9������(q��B�ˀz��l��� �2X�;ڃ�̪}�ņp��Ƞ�ٸ��:Qԫj�雑կ;�,v�,��4,��Ǜ�M�;�'gaE~�����du����p=��?u6�eR#nB�U[�+�X�Vp����	L��-������ӮA|:������qH��L5;
��>�fp��EQ6A�]�|:���R��@�/d��o�3���s����v��[�k^��(��a�Kw?�NB��nW��H�;$���}�N�q�^�UP`˻��$ 픟��`,�pk*&1FN�h�-"4��?��T.�u^�93�ߎ0��w���WQ��V��N+�:�ZO�B-�� �a�*m�>�Tr,�(�,�W���ޓ�y�Ѓh��~NzG�&��|��,d��,�L�vPu��#�Պ�(��媟�0�;�q|^%{�ʩY�o�K�~A<�2I9(���
���N�5J?ZqB�1�Ƃ֝Py�<��np�I�s��1���T�bg)��SwՏ�
��v��<<��d4@w�M�[5�;u7��Vm�cσY�`�B�k���:�IVO�dD	�|}���Y�,9����'�E�l#֦K�hc	,��m��lZր�#���U�8؟���P�w�'+�I���"��>IOMxʟ�_~�nd�bx��6��zbQ��@>�˷�G�dXq[YH[�z����5�����������@�Ļ��+�ތ��C�β8F��r��栶c9� v]�S��
�`Yv��F���L�Y�x A?c]q/�K���R@�Mk�Bfw,ݹ���܅���M���l�>G�i���,yh�h�*��u�(.i��z��ep���@��<Y������n�S��5t�p,�f�V'���e�C�ܢHllHU�'Ѷ0�
J�C3U�vL!����U	���L����ES���Ͷ�I���	�ͯ��z��:Ԝ����_Pʐ���{����s�[)���zE�K%K���J�1I�%�u�BG0�T=|�+�Cf�D�/A�x5���o0g2I6 ��α�V�f�+>F��jU(HoX	�'�p~L2�ˈE�j����Op8S<H;�A�No��?�]-�2�㫥mB� :'T!6�U����=<k��nxBK ��CH!�F\�C�%�~�`�����D	���C��5��m.�tB5q<<�&b�aW%��ӏa�*mm~;��-���"ǇsQ=8�7"����O�i���->��S�8�k�K�\z�����n�gV��+�:�c�/x~)xI[�{)U>"ƵXedx\@K+��`ђDg0)�F��<��u��4#P����㻂ߚ<��Qb�7�4�qk���p�f�u�S�+�9Z��g�<�'jZ?-M���+��{�kq�iz����!�?�
]��3�a�lF�R	t�%xߊ]�����ҏ
ODu-<��Z�A����o�ڱ��rj�F�O_�pv{��Ɗ�s�.��� `�cp�]6^"�TY�(��J>��!��R�S����Jx��(��b�q3Dě������I˗{7EB�I�&%�e�}Zs�_���0��{=N􎉯�y�/N�����Fq]�� �@5,�1����q�,G8t3�
���V-C�0��Ʋ���5J��>w'�?�F5�`�s��g�3���]q�M;|N���S��16,�Ju�c����o��#0����4��N���ٚr�s���$�ۚ����0�`�L�s�����t\�l����h�*��[��	�i��T/���b���xAv�`8��|#��������4N�(�ĸ��l�*�X?p��E��=�����;�J8��}�Ӗx��|�<�x����?��Rt-kZ�HA���\�`�|������$aŇ�ӌ�]JA�V��2�fZpd\���<:zUyM�yG:���,��	W�k�hl�+���jSp����Xj������c�F�$qП� �9��^2�oH6P�er�6��|�gi�du��3��e����.����c�x;`�L��g:�����QuC�  ����jKt�����/�J����Q��2�V<_��p�K��J�� -�K/x��U�t/�r���5���ę������L���K�����>�L��&�FM��=�x�t8Mri�����x�
*��i�n�3?��I��LXR���~yd��J	�wu}\��
�;־]��)��R��	k�3Y�4�����ז4'��왔��*Q�LdF˽�S���A����Yx�y��H+Z���?�̍���i�h�y �UM�7򕯬p�%��YJ�i۫d����=�|�#��*8T�-�T�����(�V:??-9��\��L����D���� 0�1x���Ҿ��!�V))'>d�k�q/͕�l'�f� _��/v���V!�z�M.�9����"D ��I���D�e��No�O>Vo��t���!gG�E��^+v�Ȍ�:�k�7��6E��&%��`a�ѝ� �K���l������%����A$=+}4~uȆ������N���U��!�¹&�h�i���ؙc�˸\�!&��&���.����o����]��$�C�8�#X{��I�$>�Cx75�DJ@����F���aQ%�����';Ga7��FգG.K/>l"j�n'�v�΃��x���	����@�sF��K�
%�e�{����ś��"����Z�`����2�W$��
K����W���]ٳ�J];�	�������#��'�*.�Z��z@)/�M�l�)�b��\�ǳ��PX�iuA�t�K6k�HȨ����P�h�����0j�ܔʐޔ2�9��;"�B㚿M<���8��uv�yL� ��v�j�=�0�%"̞�Q0z*�ȉ{�[W�e̥��!s3g���F��LTH��l�o�kl�7��m$kr� Z�H3�gFt�5F�Z�z2��n�6ν�.���i񅸟����2��e��܀��������a3"��[z��bv�`�@�[���L���������_�}&��X�I���y��b��'ׂ�e�?|!�-/�*�V+������X�p,�9UGso/�{�?ـ�;����~��30�j�B�	wV\6�	�T:~���d���	LO���Ѓ9d]���������M�wfG�!�
�S��3{���`��k�QQ��y�9F���+�S+�`�]��a~A�;=�ߋ�3��w�g7�A�6�n%F1��?�d@ ڻ���c)B�󌃢�7����_R֎�{��c�\ S=�!cXAQz~����XU�8%�W)�26L�2s�s�h��e�q�dT�՗���r��g��
�ujZo5W��ߋ�C4���=�A�$����8n-�F��}~�����}�ŗ�J�fe�
9�.���zz��KY�[���eK �ɝ��q,��F�^�����ĕh���kb���L�w| ��I �H@z�u�e�aϸF�;[	h|Ls����/�£�l�] 6-/��w~wptО@�3���1�=�%$#&4��<N���4��̅d���W�x�@���W�7�!?��-����l`n-�A9�����y�q�e&!��.Ɖ=p�N�~�4�z��3��!p�7�3�99�ߺ���V��/x�Q�̟�e�XF5�,�ɵ��[�;'�z���)c�8 ���/�yx����f�6'|��؆�K�~tI����^��S:���$�l�t-^W�@��.�������c?C�9��̃��"F�h�KĂ�+Ms������"�2�r��va��gu� �����.���iQ͋�fM�n�
4s�enTJ�?�2���	&�A���ô �����6�GCX�������xM��;YWVN�˫m�;�U��y�eapa�
�dr��ۡ��ݷ�4��ƚ�ER�L�/Xf�뾧��c���Qr�d뫦s*�rn�r-~'��a����x_��R.�X._lɺ�u�&7����0����~��Aw8��>ץ>�r|)��Ф*�fU�Jv)���etb1�;�܇����P=jD)�vG�����#���,��X��/��苈��g	
��:ɤQ�'�6��51~9�ucrg������y�Tg{��߸]���?����ݬ�˜6���a�0W��7״%��q��k"��i�����+L#$���P��W����Gp/��N5�����۫y�����j�"�m^=���N�Hf.nI9������\G���j,s�5���cVw�$0��,�2v���Ϡ,��O��H�ۅLoď��L�#���&*Be�����QzjZ��d�?��
sھ:>�ZN���������HL��N���8�%��l ��Hq��֠����E�,_��4:�?Я��h�F<c�/s�j7��7�Ӛ�Y�C/����fE��p�_��6":���G&,0T5��S��ڣd'7��LPJ	�,����Lj��=Y]1���v���[��- ���8�����|���V�JZ�����-*�F_Çq�6�����4L�z��z���L����	+�δ�	�Vg�����#-���<�����YB@0�����ph��W�:�de��{�g _XG��9��^;nY7�����6������e"��e����rZ��l�!n��^��&�Y��ZS�OX)�L:"�.���D]���وGGs�Ai�"{��_��Gc@�uM��Zވ����|��Ȯ��C;���_	D�1�P�T��פ����D&�_��=�V��Z�Rk�=��ӂ�䋚T�D1e{@ѧ�̩�%)
�8B��}��һۭ���C�\\��\e��Se&B>��x����N���*�8�#@�Z������߸1�f�%�u��Tb)�=	dX�0E@�����F������Qs�v�nu�f�����1��[j��S[�eS�\����{�1 �uM�B�]~�?��.�x&\o����,�����B�Ea��²�T��s(���p���&�Ȣ�����4�ބ��4�F��UI#��j�My⊟�ntq����X�r����d��Ŷ��T�W����R��v���w(�&p�O4��U���Do�Y4Y��{��Y?y�g�F�X���B\��o��U������؁�+?-��m�6D��ve�`nF�o�}�8��MFI
�N��&C�5ӯi�=sŝ�HD &��2���_6��8��-��lҋ���*�#��y!L�t��F����K�\��,�CNQ�1���euPG֗e�'czP��R���P~锂S&�\�k?��P�bYR��_��o�t&�C� ^W�{Qv9t(2xi��.M��}�b7��j������N�P�af���W8X^�-$*��#��ޭ8ឋu�ۜ0,E���v'���æ�k�l��$��ȯcN�٭��ѐ�p��Y�ͶU&�]5�y!���y�+�	�{zOU!^��SƳG	w�Gi/�T���4dދ;lcȹ�֔�i9}��B쿶N�j�� K=i���Niw*0�U���v�Ѯ�����˙��Mv#čZ�0H��#�`icMV"�HzF�� c��8-�ZS��$���l�ݏhW�X�DE�~�N"
�f���v����;���	)W>4,�7���MmW�]���ˠ���0V�՞�e��>���T��8�$g�2��~:�P�&n��C����Z/�B�7��bu�(N�w����g/��թ�}D����J��t��ϴ$�9fF�# X��q�@ok�iV���I�j\j0�Ð�D;�%�U���n���] TPQ�W����w�.�� ��ւ�I�m}<�x��f�4�z/��rt�2�B��[����/��&2��e�.��5�R�+
0��u�2�.N)�@��Z 2@w�;y?�Ǣ�x��v�Z�+��LX���wu����2���?�<���Jy>��bYrN.�5\�6u5�Ʀ
�"י���~b����,�hBa��}�Mg���&р���;O��`�~z��r�/��g;���J�`6�_�����2���Y>؄}�Fm����_�W�z[� =���p�ޱ��9B2�#i>�Ԏ�p�O�9���[ɋ7YWE�y��?�R�Qį�JM!Q�ȣ��\қ�!��?y�_a&?����x��`.zJ�uX&�ֽ`�LQ���+S+�͙�$n^b[������k �ﮟ)�1�eh��3��z�(�Rň"yY�Oύ�[h�r�5�*tS;-��d�7dt7FXB�F䳎cR��q8n����V���(�!���h;�]=7���[�4�Ec:��g;`�YU�4�;�L3t�M��� ��|�Z��8 �p\��
wY7��z1%�ԶH7�j8�IS����K"���pZG��Q�w�d1�`�q��{X
�ʀ$ĭ�3M�D9:
-��ڛ>l�!�LB�K�Y��M��k�Ǒ��R�nG1D�4"c�T�#M��{�{��S*�g&#�����Oqx�/��<x��c^W��4ƿ2�j�'to�n� ш
��f.�Y� 1����	����vw��薸^�������0�P�RU.9f���� p7��:Av�K	xB�"k���'Bu�.ܶ5�B@�!"3$<�Z�*�׊ ��A�j7m1�5�Àh����3�����'ݿge���a����loF��6y�{�n�E���q�hn�9�f���|S�\�(�i��2�c�ͬ|9�ɥU4[�|�f2�5�"5��V�-��M�]
hs�4����Hq�N�)����"���O!3�	�vM��ҩ����4�i��=8��g�hvJxT	^,� ��L�bIL�W����q�ٜ|�
&$j�6�bw��,?�ôB}���p�ӕ��1Ӏcp ��^�1g����S��/���e�o~bZ���C&�+��i��S���N;�<H�5T�"���q#p�%�	��$y��f��i�S$yyO&۽P��V��������˟�d�}+�:�|z͘IDs��U@�6u���E��h�taK8�K:xD!Έ/��Oh���ܴ���xROKCs�{��M��w��}���+z�5�
�FD�����:�%:�7��Rfb&W�鱧gN���TL8�~FlY�����~�X����U�'�� U��I�@��ץ�]�;4G�R�|�@BB�n�쭇��ʳoE,a5���s;��9Xu���DK|u��ca"m'(����y�>�_�_��ϊK�<��	@�bO��ّO�`�R���ʼ}.t��"���Yt�=�J�@���U`rq�*����)�B������U����9�p�I�PP	H��iӑ������:�Z<+8���ȼ��E�ֽ��2�4Bc�°Ã��%�X�H9W��-nȲ;l�[osOrTX�T�X:O�,�J�muFƺq����#�а��@�Q���m�jHF�e �jKs8O=�H �,�|�����7R���*ъ��P4�@��u�<����0Ʀ�>U�������3:�NS���?���eg"x�e���h�$(Ncc/,+�^\����1��`�޲�o�i���1ޝ}���=��`�1}*�x]v�u�/�EK1��Q@�Uw���I�x��PT��Xŝ���9��~Q-�՟/��y�i�9���0G�&bq��v�������ݡ�Ù�YS�"Jl8�n�e��r�e
2ÏX ���/ � H�g��vA���/����\�%mbH�q���8qB�H�9i��&�@��F�Hf��5�2|��|��Gr:
�����w�3ݞ}��q�`�PD��Q�*5
���-ԯ;����:��Mm$�7����O&5��}©oM�JPK?��ȠR�G'�Z!>���k:��
��VDcO����S��`�aV3��L�Zq�ᮀ�cr�OI_
O,����4�-�����,E�^��������.u�!!W�f
����Jk�@.�RM���~0��6�E4����#P;[��Hd襓���ac:>%�Y=+G�6�F���5��&���`��`�FC`��ykn`���a]q5�K�����b��,_�Ê�e.@��n��R�~���O���u9�J�s�;i��N�pQ������9�*��Vg߱҉���p���P�K͐ɉ��9�I41eA��s��8�;I�C�v�6T�|�8�.I"#Z��0]=�dM�SC�)tz��l�����BP�#zb ���+�FZ��h-�H	w���8��$��)��D�G�^~�e{�I��Vᢊ���C.��c��9�|ܤ�(j��.�t谪8e�]ׁ���K+�OR���K�lgBHզX�M��"E���mKS�]������ԇߺFV�*1��	|K	��4�!f}M�&���?iǟ']��y.��E*DP��|Z� �f��ı{�;&�lޏ+�O��3I]9	q��$�5��T�`z<�����e�vT�i�,*�k�r��S��?h.�0\�����/Eg#b��5����#ޏ	����A���q�A��@�r�E�VF���1�	��A���%�#�`�H�..�ZM���m0 m��8-hnZǦX��FM�Ͻ��z�s���E_h{����aW��2�z�P5˅k���^泽جͿ��C�/]�^4F=�'����P[u5Jqj╬IN���	Y'\nꝱ,�WU�GS�I�Ķ����=�L�1�#�V	m�����b�%�#�^NK�GNt����̋����`����MZ.*{��Z�{�K����ٝ�I�w��1�I�1�uT%{�B9��<#��$Xuq�9l�vC1� ��?ۧ����]K"� fh'��뚴��N�w#���9<���W��O���7"{���t�Hpf��J�[��_V�#�"�Su)�l^tfn�����#04sip����bC+N���\�<��s?�ְ�]�W��P�t����x�p�,�@�&�^y���s�(1XF8�2~�
i����p���%V��^qh����^����k$��nj�5��B0����$#�7��AO!���o���.~�$`�RD3O3�^�:M�~�SY{�����MGy����b��@b�W�7CC|k�x����Z�`2g��C�Z�ʊgЇ�x����օ����I�u�m��qg�,�d?-���Z	]�^��KQ'���]��Apc� \X�T�����!:u	�j� ��3ج����(>��H�)�����P���g.xN�%w�	���0���H�sY'q�x#.�Ao����I9�>\����x8����.NPᐄ�'�Bb�0��� �x��T���~���Fo��R{���/\5�֚#~��s�It�i�-E�A?cP.�S�ߡ���J�]�d�?���-�	WeC�%��B���f��R��c_��O��Y>C-1��8�R�,��[�S�&O��c�����J8)�qA�6�rTK�������5�(;���A�sy�#�e����7�~B��oi�u+J���/p�V�H7���a�UTX�%���co��Hp�Dh���J�������`:aT�+&[^���QCt����r"��lS����sǲ���v�j�8�P[T��Z��?��R;IZ19RfL��4U3�>I�| ya�+�>.��(ƥ�<'ĵI������N�	�dW����6l�L����C�T�/���u�1��x�3�{R�	yVqS��IF��C�!���σB�� �0��Dþ��wk�%���p�e}��^;-�V45���gp�.���߀n�i����z*'EPLՔaz��m���,ŝ��%�~�5��xb29M�Of�̡n���XB���1y*JZ����{��L����#8�ď�FB�z��Z*�)�0�����-�d�d����������b8�:��_��~�~��/~�_.&�� ��r��0"�A;�O�eZzha�4���G��M�nk9��w�L�90U�N�hEp&p1��=�]��<ˠ�j;�KE�����e[ό�G0�D#`C'�S$*�=3�PK��s��&|na��>�8NX��°^C�2N%y6Cy�DL�6BZD&hD�v`߿!��B�z.�ȏ4�]�!S��8�Q����Ǒ��Ѩ&��4�}b�"�E+ħ��ZCP��m0�1'/�|��b63�$} ˏx0�n�-���D�!�I���f���F��1�ў;�'Ic���TJ,����%��"���$|I~X���Z5���3F	{�Q:�D�����B��iS��B;)^�\�C��P�]����G	��E#�	��E�Js+��鴇λ�b��xH���b��z�z���+�����\�x���H���z~fB�fX.B1#V�C]YV�#�l�����a�ܰ�t�v/�	<���)� ���%U��W���;
)�؊�0D)&/���S���I#��H�s�"��R˳�ɬ(�^ ���@����&�+�k4PK<�D���{�r�I�l�*h�ǽ�:�!�[�d��ӛ�2���2ep>�h�5}! �Q��)�U�<3�T�������A��R�z_�Y���ҳ�q������m�<�x�D��f�Ȫ����%�~I x��y��}��� Kz�2�<��4���a�����0K��� { ����h�ާ��.��u�36��](��c�K-��W5\�/4Z�f.z���ӢOש�v,t�'nt�&��ͮO�o�B�����`�޻.�}8��uQ���!�`{��Dۋ���l�D.,�3'.����������"�'/|y���yJk�
g�z��L�s���~���)g��U~ڟ7?�G��+{gN�wI�rq-_q��?53�(�f#�<���;�5�(d0е����mi]�t��;��֐9��k�P��A��X
2���d#gY^V�g+;"�3/�9`!�*�(:��&��E{^[f&E ϧ������Xb\�]2�,�޶i�lVDk�8��+~��j.��ҷp�
�}):�C�~h����l�]���� vzgτ�&<a^IY#��i
�N���yt����'�?��q�P�Z�v������!�EfP�����Y��P�F<�)�PZ硯�u�#����
�����1��3��YV����Gծ��b5��Eb���tg�w�L�CO�
�df1s��^�/sj�:�˶���L3��w?d��_�{'0VAy%B�=P���8�5���xH��lhĢ�V�R�v�>h�%Vw�7�n�Sq6����@dc�::]�l�H�yƣ�ʶ?�h X��f�l6i?PP�r] ���F�i>V���wCxO���Oaa���c��,VD��s0���3YǁAf�*S���}9JP���H�ZL�D_�M�~�m�!���e��������Q�Ǖ��Sv�o��8�58pּ�[���k��9���_�P�F~v��; �۹f��$�`�T��&y�U}fѤD��@�����qa�)_��:�+b�_��G�L�,[5(��"�R��r�jY=g�S��3�l (�>t�T����48����g`Ue�G�k ���\���A�	�j�!����Q�|x��6������@�#�?�U�2��c���WYɦq�f���;�v�V�hDl���Вr�R�v���r[�>���N���?�c����FV�a�آ\���Zq��P����v��7��k�?N�ncىSYf-C�����*ȯ�mՉ�6P�Z�h��Ű&y��{5��;���T4Ƈ�b���o��֫�lZ&����:�>NZ1z������44��,~���*u�l�q3�"]�T��/�o���� ��H�5�4��3�W�هp���S)�l��)՛<X{�qwFQ,|.�G���\�1�h7�/ģ�>�C>�hbZ��	�Mk�J�����zm��̠��S���]�3����}lk�)Ux����R4؜�Ny�͛�����L��a?�͓��v!����Tc�$rglP���V�;��qu�&��x���;e��Ӥ�X汻�؍�ot�d�s�o]��*�m\|DP��vNm��	Iq"�G�_�~�̌j�9`R�M}$1�'�N�t�5|rR����~�����o�,Pu%>�}������I.T�r�ᕥ�'V@�UoL�?@�<��SlSm�X�R��TK�Hk�*6QMq��j\?.+�PX$|�d��\��_�b&��_�T��D�[�3���C�㧮i�l#�%u�m�@Ū6�yD,w��eWGs�6�i�����~ni`8�>��UC}�=❻��"4US�&1o�Ξs��ZÉ�}��1sA��<=4'x�)���8�w�f���
s��R������Tג��)��}�MQ ؟��;H���θGP�����2�����U�i��!��Re��H���B�R��鬸g��mH(LH�Ţ�i�b��2��v�)�|`���ABi,�4�������ld:���MԎ���]��&���ZE�K<��h��8�@��>c>����H>����m�M��x��^�/-�wP��e�O��|�~��KY�'�j@��q5��7��2�V���˙$f���ʿ5,Y��A@�PM�:;��[J*��ulr5�o}	s���C�v�U���Z3o�ڰLrt�Wΐ����s7U�/ ������ ��4���uJ�o`?�A:��k6��]����ܟ)�IGڷ���a�N!ʇ��<�L~�NS9��.	q?���ƂӚt�������5�!Ja�u�{\�**�ŭ���>F�g��N]q��x�LsW
oMnmo}Jk}Qk���Y}�|",���{O��d���[�_,�;���6��x�M4����S�F�7�e[�ʛa�n.:3��~�(��|�M�v�\L6h�������e��ٕwS������)�UA��`�9Dׅ٪F�	5(���mw���-Ê-��g"��,�s5\*��0�_�H��3�k �3�I_�❋�qmT�rbc7��WW����z*c4=�)��F T�"�[��"��-'��b$�CУ�Z zF�0��J36�eR����R���X-���n�Af�zb�C�3>�ɑ�5�p��2�\�C��ɋ�o{ن@�}Djr$��.�	R4��d�-��4��aj�xD��W<���?'��S

W����X�ٹ˜J\��;���#ٿχI�V�X��׷Đ�������a��:ah{�d|�������u+9w-c*�����>	�L���vj  �u��NعaT͛��=��L{��i?�5vڈ�xR��_�a�>��Q���y\8O։X�r�&�C@>�ūq
�N&h��8g}�1��uG�ۺWp������;p�E+Ք>�=f�f�_�ޢ5�#A�.�و[]E��]:{�7j�_��/}�K�6	���kOp���N'���T�����~n( �k4A��Yh�*�_z�����u�Pin�A�^�(ʫ�C_���A�I�\��� Z3�����D͒��Ws|.�1$ó�o����$I�}r��T��}m9����Ȧ0-�+*��@�eΤk�x���p��.�Mū܄�NN�|i�e-�[ SKX��ɻ%��A|R���4d��R�����]�no�}�M�>mA�g����dE0����@ tzf|����:"�%a<D�:W�FU�7H���C���z�����!�h����}��C:��btz��YN�h��oٯ��{>��8�\`���lES�n����T.hM��+������ɪ�ɿ�a�v�bˀ&pV�}&�|���c<Gi��oB־�_�t���}��������q�����0$�V~��B{��
�zyB�_̜���b�o2u���	Z'WU4ķ89��+�X���8�"���(�~�����Ŷ:�`��
r�����F���T��f1-x�g�C�d�uEPho&�Gӂ����2g�����'įbwy�p��1�Gq�I��0]����<Pf�.t�"�G���*�6��h�TJZB�l �"iB�\0�,��)�3�)�ho]��&�1������r�P�˻�->(@Z�v%�������!1�P���^=9) -'���!V�J�󚖰-��"�!���M���H��6	��m��U�kCt�6�P����()X�v��$�m?Z��=����aa	�-�e���%�&ބ;m"��6���	
����]���e�5QJ'=��&~~e���6<F�����$���KCБs���p��u�Ә�2�亄�{0A�4]�Rp�#���]��n�d�|+. Ć�(�M���f�C�~(�/d�<Jx0�ۥcA�13���%�FE�d	:�nD�U=�k���o�u�t�V]b g�KR�Za����J;�g9����r���㑰> ъP�o$�#O�p�����3᭷9m\!�6��WÛj�Yn(�+uǫQ�64T��hCq��>ĘŌBEv�	ǀ�2\��đ�f���L��T<� W������ҭ�)l��{v8�3���Y�2��P���9�$~���}>��pC8�g �ΩӢ�˪ky1 �L;�n���3Y��CSɴ�W��(7�; D�q5s�(1�8 E�b#�[�߉�b
1!�m �E`�z�unn4���wMA�4}�����A}}���2���pLQ)K�.k�Z!e
0YTm5�T�\�a�4�|53�����2N�%O=R�N�[���d���M}�lu����\ hY�'1���.ޮ�CՅp@�F�ACҠ��c*=�x>�ŇM��C��(��W5S���ʔB��k���h��G��[�~���A�NO��C�L���uzE{)�%�|�`��a�l��.�2�@���>ng}�yCR=*�y�fC��1un��׈s����}��G�z�
��a&�a��C�|�S=�N�M捻�&?��x�aAk&2";���E;ԲrJuq�P�֮R���j�KΜb�r7��ƾ�=��&K���rJ�)�Yj��M�KH.���Q2����ΉO�:+���&�L�7yxPС�;���;{�twY�n����^s��B�nf�>��ܮ�����n�h���8���m�����P[��.�[�`�U��?�/�R�k5�b��R�����@�R��{B,�sW��9�~J���Û���Ճ%��H�*�3 ��9n���YG~�\�n���j��;u�uP?>E�+?�V�Y��&0Q\PhlZ��1��l޿�S�P�:oBu�����鲌B�_���Ja�D���C�^o����Py� ����3\�y��Ŝ�"R��3:>*��� |����X����R��Duy�:2
�����($*A(;Nh���������Cr��#��x���K�SMH;2S㬉��Z���T�S���K���g|qjN�Bn�� ��T2i�[Sk|t����b����U.�t�Sd������p�ɚ�B⋓��S%6��ڶƞ&��ZE9Gb�rt�%�û ;a蝱K�!�� c� �{$c�p�9��i(Z�mIK�G�I�JXz�UX�~l��e��IJ�r�����{y�Ȟ�}a�����h�)�8�d<��B jk��h5v�
(�-��Vx�����W��D�'=��׸������/�����I�M�?W��a�L�����覮ք���R�q�R��]��מ�5��Dh8v��Z,�}�-����E�)X��������̊���<g����!w�đ����R�T �&�]}l��b3��p�Cg{��k�{��4�ν�{�Jq�ZL�~�k�14`�*�X<9��M� ؠ'���ͬ��`~ѐ ��BN��I�V�;�XnO4~��z���X�!N�.x[���:���$ǫ�Y�Y�:��= B���d�#�.[ɀ�n��,���<��q�wdr@���]|�3�
�r�����v�9��j�\�	*�EgV���8[K]F�ˡEv��wnn���^�
�Ē���W����N�W��:.�J���}�t��i\)��I��ٲd�8����#�6�cxJ1x�H�6�jP�I��ֶ�D2"(��0�L������ݐ٣��Y|���4����W!H��Ħxm����#�֚��;�u�v�����CD��h5{ΞG�x�~��s��'%�﬒��b���*A�5C�/���2A�gk��p�������U��^�W�������̉N�]e¨���1 ut��80iV�\�������`v	?�k�'�N0�/����ɛ:�3����Y����3!~x��{�١�k2}�w���[��H��a#��Ղ{N�2G�7[-�+�}Z<\"4�O�-m*q=���In8��`a�&�w�BA����Ny���(���H��D*�h��囹�5�lR�}C�*At *��9�G��v�$��IA�Nb%�L� �Y��t�M�j;�k�� Ch'�lA��Sz�z�ajO]t��!���AńP`!�ѭ�R�-����,�;w�V�|Ծ��: �a\Sțs���_�^�#`[�M�73!w��Q ,���9"�Q� �ut�V�Ʌ����j/Pc�E�}�)�*_m���\*Z'.��J�,�-LU��	��B}S]e���r�ëC06NW?�TQ`�/"3v/�����:�f�٨+M�(A�L{�y���?�42H�UP�OPB��x����%��gk���&��k>��ڂBhB�!3[�%�@�u�R��*�'��.����x��Q� ��˯<P���!�?VFV9�I��-3H�a��j���H�[�N���/<;����ڔ�%��F��X&Gu��.h�O��E�*���b��/�!� ��q{?�� ��Z���&.���3��M�K�9: W0{d�5��c�Ы�G�p�VV� w����&#�����5���Z�=i�E;nK.�Q놱#i(�����=�[:\W!O���9���t�͈��:��ID�06��(ܮL���^?am��^_���ؿ]g����hA��?�����`z����~�	�~�aA̛��;�X�8E(aKP���������ȩArQ�"z�H`a�~@T !p+�:����79z��A6\��eN��˶F�w�����\�A��=Z�eX���-�)��
С���W��w�To���7V$����'C]A.�N��4?�l�v�!�oi(��A 	�������v�q65�*�Ԥ�(��t>.�-b�鰤v'7��g�J*��^pΧcn|�G�6d���Ym&NLE�[��yg�D��:V�7׎�6��~X��w`rc�{~���޻Mɖv�v �f���Ϣ��=�OasU�:��Yvpqj'�J �.*�8u��e�,N�9�P},a)���-�&�B�F�R﯉}~�lBb��y�&yJ��¨vIw�őR��`��I�g�]�؄>�f�W��8H�8��)|P��.�Z:G_5Lc^IT���|���;T��xǶ����v�1|[���@�����E~wgE�$cś��Z��n�y�up��s;Bg�I��"S�YeiZ%�~.�ɦ���}���g��Sv���]���댿4M��w�bo�z;w�3�]D	�m�X�@$�*ڋBO%|�����&^5�`$R"7.�c��J�R�Jl���c� ���;ˆ9R������F��n��,������:}<��Y7Y�h��v��S��JCg���E�����H�d5�sB�<	�Ī�~5?�P=���X>�t!g���+���U�ʚHz�m1Ep�x�/34�~l������{o�����-Z���
 "W�ȳ'(��a��jp��C��P��X�7>�V�i�7��+)�O����6=��5�A��B�k������2�R��\}w+�24=j����Z���0>�R�f����i*�����3�oܷ����] ��WptT~����Q��rX$;�<�	��l�[|8mǵ� ���>�S�.4��N5Ȓ�j�S���,���s�~�gh1�&�FZi����q��]���]�w��<�B\�:w�p'�;�,�����*�f]�%=�
����d%�8��۲] ���k��2�Ll�i)-P#����H6���(�=���B"S��!��h�c���Hf��&(x�J���h�a�K��.��>��Ѫ�D/N8�C��r��J"��H*��)@l���`%�E��O�qwJ���_;�Tl>s؅M��݊Z/vs�1U��9�8����NE`���]rG�?��jI(1r�ǃ� �8�P�O󥞌���(�Ie3[�JP�&���S�	 ����&�$1(�����������}��-\���V1�@�fv�{����vk�7K�!�+~6�6t�ϭg8�sPUOm����"b�/ ]��<��(�枬�䛛����w>��6"1��|F`ۿ�>��'���& +�oݽ����W&���t�/���;�'������ߐ"����,�k�`�Q{3�:�bʸ��v�g��p˞)�!a��[�<>�?��H�OA���P�zC]p�ψ��#�	�*�k�.y��mG��L,ZY����I^�"D�̯H�~�eж���3s�Sf�+�����6���	�W��__��l����#Aq�}Q������r�Hȝ��M�f�����i��d�2�l�5D��%Cʊ�
�a��f�/��9�PX���	��W�ݬ~���[�j�"�>����d�\@����~���U�{n�hf�Z��N�R��}�����:f�]���1�$^^�ѹ�;YJE��ۍ$`�S���6DI\#(�榢���J�s���!�EZΉ>eY��I��D L*g��*�q�k�O��9y��!9�w���J���������'yD��ț��X��8s�l��CE'����Gw��q��ԤCP�Ή1*��!U�����߆/m#t�+�0��O�*��u&Q�%T�@S�]9U�2e땙Ĭo�D�0�����Y5}���)ͳJ�É�Ǧ����늆w�)��n<�W�,�y�ߓ�J���݄c��D��3�:�I�����s��?��*�&̲Fm�����|+��U�`*]x�#I��c�Ԉz�?��d%�tP��,�]nP���o�5����촃Iy�O'�l �m���|��&�:�re����6P^c��P8U�^�D�$�,
�)�>� �����	�ŉҽ@�R��$:/w��%L?{�>1�+��N�U݌�2r��6x���6��
=H�����e�7���T{(�n����Y�w�)e]6Cڋ�L�`al9�ىI@2�O�lD�.��c=@���C�=^ӓr9p���]ތ#t�<���h���36y��*m���b�Ho<>�G�Y�ȇb��6��E�SQO=14�o��b\�(d���EŢ����(�5�'Q�׺�_�u��9�}� ����8���f?�6���=[Ce��b�0J%�/�|y�f;,�#�W|٫6�mPo��=��[�g�fv���KmD���c�IN�R�QEj�q�مaJ٣�M��HHY�� �d��_�|֑RnĄ)������d��D�/gM.vf	�0�0���r����PZ�P���V$���I�儹�-���z>O���%��k�2��}�	��R=5b����Y��{���E���S�h_��N*=l�+35���_h�`qPήXg�idF���_QF��[�ܜ0'9��.RF�L��9�ӓ��J��,2	�x���3k���6��¢���C��Ou:� �������Ձ0x�W2>UZ/���4���%Q:�sZ�Ǆ��	�
-�n�2�5Ƿ��!�E�.CF+�(W��5{�O�!��k�L���?�w�1��.�����P���W֋d(�e:*�������q�o��`EZ�`~���sS�x(���|T�	9������׽����?�X���VԈ9��*Y]�i�ʑ0Xr6�^փ'}ˀ�#C���#v�&澉x��A_�����u��Em�(ᇲ�vTC	�H`��z���&�}A0��{�PÜ힬AW?FzÖK���:���vay�|�`0�p���;a�Bj��v%x�E¼H� I�\3�?z�n����(��3rM�������ԏ��2�~J��R�<�AQ���K��j��6���B' �DT������]61~8�]Y�`Û��Ք��[��,¬�&���F�ItѠN����4���/
�%���x&Ia�e7���`�����rf_nq����u�;�f�p1|�RBO+��moW�����/ȧu^����ǚ������62Ws/�GӮY%�hdeU���T/�S{���]����D�b{*�J8��M����d8�fE����ƃ�٥w� �˛C2^�d!��W�� ��h]�����D�4�JR����Ą�6�T�2#(�L2���z.�X*,~&=(]�w�e�R��� ����G�%��,�����y6�6�B��f���5Ɇ�(�ώU�q�I�t_��A�K��{U���ߴ��+a�/������e�9 �P��)�h.*���U������2]xc��[6���G�T\�3����,�F���/&�����A��D�<�
�˛�W����� 6��b��ށ��� �/�1S�7�x��v8��X9�d��["�;#��NRl��5�i�vA����U���,�9�'|���j�-W�s�R�V	N�Z��� av9�(�AAU��E�,�@���t�׶�7n2'�;EЁ%/ox]��6N��_uը�
s�SH��`�+/i��du�!_ᘬ�AR�f���βɷc'�CL��2s
Rq�;]o��1.7�G��s�����]��wspq�vo9L�F;�9�"*\����?0zͪF9��Qō��������)"��OO;Lz��:�]�W�(�T��UCޒ��bG��}X����Ő8
D)r�|!]e�b�3�m�e@>A����l���FpV�&����Ȱ�i� W��O�Wȃǘ�[��5x�����b	2�G�v����e���v����klcw���^� My�&b�ۑ~��\%�L�[��e�O���E����{ȃ�i �����c>�y����M��Tv)�4P ��J,N�a���}W�l�oX����}܁�`c���oB�h>��m/�r�I�q�1����|�z_��,�_	WF�c�6�U�Y�a�,���Vs�xK�r�#�+mv^���?2�>�*�납y�n7���kJXP���2b�Z��c`ѭ�r.*��b"&�|,"����a����r�v��3X� 9�"i�,~�U<���&��o�s��.íVz~��3���w��$A3�8L��R�҇�<֒J/(Ȣ�jC\�d�:�kh��۔�āe}�,ޣ��P�i����d!�u�W��I齦����F3�X��V��V�~�3Zӫ�f�K)�j2���hNE���
� -sf�zi���]�8�2�xA�䘽�9�ʳҟ�t���&���UQ�饊����!���/n��Bo��H0q�(�]�l��:�Ћ�4T�e�ns�׬9���&E �ʜ�Ax0�_�y���bu�9�s�S(o���H;�)ðl���n���G-豃_�y�H��z�"����~��h-l��C�(��;J���ov�yGdfG*ً�[M�:���o�aι��A�~h�K���a���*���h��RSz٬��������q�D"� �bkZ����l�LRc�Ѻ䧜�R� ��	򩙔
��}�G_9�}�q)�H�@��֍��@ģ���`�Ayyۥ�_
`c�W��*���/�(�<��L�@�t�τ���*������5ŋ@�OR򱿞��`��7�9����أ^��1���Z�_��M'8_���U6Ec��eEk6����	�[���)qex^�7�')�F���b�'�p�xB�"B�/��_Aª�<A�����z���Y�? t���e�G-tL��H������.��D�4�� oe%KV�o?����bs��D�%X'�h/d9 �������a�X��չM68�:+��Z�XN��.v��� �]u8�λ�[�(4����f�ɼ	KN��845��zR���)Y���Foe�,!.Pu���@���焵���j��62�:֊fd��󸗜�UJ�U��'yH�#$��ұT� =X���@�(B�/�c%�k��|x_uM}K,�1z�g鸃v7�]���m���X�0���u�c�^�a��p� �$�m�/�r �:P^�ʈx��h}s�<*���&W�:�V�������!"-i��G��<aȖ(�{4�~B�fˮ]���)�(��]��	�	;�LD�w�V�ai��N�Ȱ
��j%��������FW<�_�4���E`�c�
�T����}��*�g����k.�����fb���e�~�K���w�� H�e�͕;��,�j��C��ˡ���7o��GC<m��|���~\�+Q�И}����ň�|OA4!��8�_n��ﹳ[`�+��2��桢Xb���`�/��g`��3�&��L�X;��q����8|j�F�w`l�����{�[)�i��7�=��qz�U��ޱ���b�1e=�+����j�{�8��E\OC%8��9�i�I_/�s( �rl[J�_�{�:%�<��]͉�d��\8Z���eI���ݝ{�f���� �Hy�G���������K.��u��1d�>�y˓>�Ź�iۣ5�R_}���YvU ���S�M
Y]2�ci�˖VXoe�j ���<'�;9|2C0�.�g��]��	 ���M	T�'���Ð{B�����|�b�>Ѽ%z���ќ��m�%�bt��fL����r�Qa����;4<��4� ��=�J�hQF�kP�+�$��3rj�*�:ʄ�_s�D�"'�{~_ys�!�IF����P@�N���ʰ��c�o�0� R��U��9�m�w�N� QY��o�f,�?K_&��Y���əbӬ�	� �9{ �s���U���	4FI@�Ԉ����ߊ���My�b&!��U�E�%�F�xc���h6��bm�]"�xċ��/��HJ��g�_�f���Ԍ�ɇt�`�.��UekKTTv�g���鞜�5'6�S���R�ʖU��%��F*��ՠ�ij?�ө�e�U�O��Ճ��|g���5.�vi�>��Kdv.Mn�n�]1R/K�#�����
�㐆��.0�����?{Ə*Ϭ'�~��T�@�F�>��� W�.����K��Bı��҃7Y� 9^���V�R ,����I�K�f����vI�s��1Ӯ�Wʏc+���4~H.;���9�[�v�h�>�c�KC	��DG�D4�'S�K�.�8joZ�d�8�񐆬V�<�p �h%kc��nk��UQ�H�2��
���w�����>�����BSn�u�Y�ϧ_�Kx�v^{������&�F��e�Yi7���gК�B�G���,Ty�Ss_�_4�����&A�M��Z<>�gk0�,��R��?Z�м����a-��~��
Y,��]|,N���n�J	�?%����i<�Gᰘ�a�~L��=�.z�
�<l���ؖ%�E�C�P"���*o8�n�A����hL�����%Vd�q�~w9N�XO�X��{��ƧaۼRmS�3�;H�]5F��"pX�j�n��W�p�M>&��?Ē�P;�a9p���`_��{VU�+4�~p���/�e��C���I�^A�,M��0d�a ���Tz���Rj	���ķ9��+�I|i����`{��wQ�P�q��k�'t�2�2{=��letƸt�֣��il�9��c��j�< آN�(�����h�����!lU'o���j���G��Ѯ�3>���\<���b`�74����!Ly4�@I-��~���G���tƜ��<(�2��R7Wbg54���Y�EZ=�݇M�˨��B���,ң���Gp7��]�C FU!�JεE�"����a]h�L:����D��y���%e�-��r图|�|�l��`D��f��^��ޱ���s_�\y�@ÿ��ԲP�L��-c�d���Z}�D���1���J�J�%��
����!�M�l*���Fl��d�T=�Ox8bzd�m�c��@�p��ç�q�?{t�
�IƂ9��R���<�0�5~�UU�;'dʎu8�b�~�όF�y��n���i�?�j1fИY�O�0J�i�T�/����G��ȸ�!7
�#�==y�]c�\�)/��J�!��%�9�fq�B��Q���������(TB6��")�����z+�<m�>$��֞�j�B�h�׽�K�0��C%s(�3�Ke���C�@�T�0�9X�2@a��N\���Y�����*+�+��Xލ����dS�_��Mu�3~Y"��ˌG
������I<�l@ݠk'Ѣ��=P[L��c�[�=1����Zd��T�KI3
آ��U���o�n"
LA$�� e��E��)/%'�r6v�<�.�M(ʡ�T�*5Q<%��9x'���R9��1�^�� \/��Qq�^Dc���m����&�b�*t�J���:� �=O�<;r�@Ϯmǂ�N@��K���wA~��������k>P+�^X��N�-��`h�Ɉ���6[�"K0��3`{~��´��n:��g��$��:��F�$�����^<P�x�o� +��j_���TO��� 	�d�����L5n��b�9{�Z�Y�G·#��'�ZX������8c�W�'���Z|er)"�s+�	�$GS>(S�㴈s��d֩]����P^�=�Z��ρ/��m&�1)ɟ=�ܗdy�S���SW%,��q/q�8��a~�-D �$P-1un��?��4L����v�r8`f=��t���!"����C�us�9;|6�Y��n>����^=���[�4��������(�4�/�pٺHѡ{5��"�ɏ�b� b�"�Fr*�$��
�ٞ���se��"�u���w����ic�u0Yc����ղ��SC�J��5¹�"8���E���C�_/(��U�(�M�y$��580��߱���=�%(�n >�o�$e�/s2�
�WS3 ��Gʐ:��C-���	���8�ڥ��N�?E ��gc����%a��I���k��ʟV#��Q
��,K�y�,�wwE!p%�Yb��2]8��Rz�I�s�q�c�U��Nؙ��5�5)e�_>��x�j�� �ő銱o4�W�3��/�@�B���=�/�Q:�����z�N�]��PT��Ƶ���&]&{�4$ƸwѦ���n�xd;�A�Ix�}�m0Z۸C T����%s��y%�R�8���h>c�㼼o< :"�8z������ ��-67���n�$�9#��-��ng��wŐ/��F�7��A�s+�x9*f]Ʌ>5=����T�J�Z� ����sd� \�㺢�,�N���@I3A�ɿ�������&�s��4��� I��
lL�EQY)@/j���ȹ͇6Ճ�c��ښg�4�n�h�O��i�2�48�䦤Z�>�$ �>��u���d�X��G�6�.�5LS����H�~��i��ҟ�O4��	EyǼ,�,-K#�&�;�/������I�t}�Q��X�?!Y	��MfK]��aμ�R�����ƇD�qUB��<h�ɷ+��V�P��Ӯ %��)�9L$�X���m7D�@\�=W�%1Z��h�Z��e�aU����D��ߟ�6�WT�	��g+ߟ�a�V�=M�JkS�n�O��?����@�u��VuMY��J��g#[��������9E������N���an|['�4Dh��qG��2E��f�aS���?2o��R^F%h�[�E6s��r�/�λ�ܙ������vhY�:	���Vf?�q����&|b�F���zzG�xøQ���G�i"�?	*�����u����!ey�{��?yq&�`<� ��vZ�,k�����	f�_��su!��3���c�{@?���yt�Au���ۮ��F�$��!��D ЛXv� ���/�� +�4�bqP�?���P��s$�U|�v�p�y*J�#�㹁Q���0���]�!B��$O�E��6����1���7A޺U1q�K���}��C!�%��f:ǉ�w�5C���<*%9�ls{tR���錣���d(��*��K�Kb�5��x`��{�Y���׌�
��ht�G�u�*��p����g
�+k�A���Zra�L;�K~�����w��?\��KJ)��,�;.Z1��MX���-�Sxk����9X)�S��Cy�(8�:Ə�m_Ҁ�>ܼ{[�<7�E����XTjL�=Tϋ��{��i�x�����E�VC��l�&�y������_����WG���aX��O��ʒ����i��������L��(�y�VO�۩o�0~�qL`�D��M��!U�.|	�A[&Y$5�'��Kʖ�����X�ҁ���;G(��W�f�d{W@��?��<[H��(IR�p�_�̬N�sZ�F�6׽�33�/��0N�~5�:�}f3K�)BhZ��c��B��fw�w�$�F�{tSD1�`D����G�{!�����Wq\Vd�xW����F�t�'����ҡ��b����e�Aӛ�p�7"���I#�(�,��:O9`��~�Vn��t/�'Xj�� �ڣ��щץ��Ү���ﺘ���C�:����n`�t@N��v!�&��4�o�z_��w�p�h@ѫ��^Ԩ,�d���R_x���z�WԼ���hm#��]�|\B���2!�;�O���-������<�w�O�"/&f0�Nob�յf;�_�M�}��x
�ǩ�̡��T�s��&!����n��J���� H_�)�n"��D�=Sq�[LS����I��Z���ȴ�VC�\;�n�
l-t�~O�F7[�Pt������wy���@3�+#7���.	�_�Fl���<p���`^h]�dP�T;:��-A����1j�+V%�]䈖�b�R��������?ks٫Z8���-�H��!#2��R���C���kч�P��<��Y��H���P�(��7L��=��ؠy�*��]׽t���T��oh�G�N�e|Q���6�)��ꅩ�%���x���d�ߡ'�+�sD�_�3�vM�ᾷrI�<p8�uW�����6H �CO,J���*	u7 ��W��-<@�Ғ�_R�Z]�8Xhj��:��!�E�R�{ȳ��G7���F��b�lX�����ܤ�P��<d��+a��������0р̿:;�*\�����O�(�K�!�	2�h3R�	U�Tr���SxfY� ����9���{_��Y�"���Z������X� zݙ�ҵ<:%F������'D���"[�}��qD��kI[������^r�l{]��j���0�NV(߰��S����(�BS�^��Kg̮~;��ѕR�e3ʟ�H�H��{�<
��ތqz�Z�0^�� ���N�*��[Y��T�y/�|�Y��r���'�x��56~�J�O�j��fTE_�4SU�B�R^��:$Q��Ǳ��]<���K}����ՄpI��(�A�	�{��ըw�vV���hL�@��Ԇ�7қo��]���;Gu,}q�,�6����箚����
�EӬQ�t?s&��/��3��{Wx�u�w�����Tf��C��y��6�.��bk9!��Cb�Cq�##s�K
�����������n��/@�\�2*I��D�9��07�Ж������Z��W*S�G��;qV�c�J�y��8��í�(P��=C�9	)�V���r�Ȃ����B��pv��r$�%���`8`� G���%Һ�RҎ�m@`Y!�优����G���1䴙��,�w� ��$�PT#˰��N�Ė&~O����yL
��ܮ�}�%1b$R�C�f��3bęYS�q��#'D	�'�8?p�֛��LH�_%s����P�[��T)��qlV=�!��N�5���݂���m���@g��)7���?�^�yR�44��q��0����bٌA�X,�,��r�^�}.�R�`� ���NP�(>?�ë��/!�D�o���7;��邜xh�*��O�$����0^B�����fN H�Ӵ�Ƃ�r�М�Q�9c�L�>7�*jU��%�u�˜3�2�7��I,���/�:����bJ���� ���=��� �*���f���~N���i�TR��O\P�΀GYt)b`� z�F��0��3�>T�G���{�)κW���ɳ�f
���}��,L��&T�ۜ@�;�BI��a��]������{73�C!hV��[��O)w]�|�����Y�,S�^������Ũy�<x�ٿ�^2t�	S�2tu�	ON��&XL�^�j���eւ{4A~��?��"���,K������>�TҎ�AJ�(���l�D���1}�kbx���|�j��$V�.+?�H�C�}�2�F�:Û�g^�R��P��ћ���o���ߐ� �����K#�E'�>�C-���&�Y���//�/9�w�=n����'`�["vT#�#gG=�b��o��m3�)󗃝����-��p���c��v�����Y�p�xDeJMg��  ����67��z��/ �\��@�r��7y)CO���&wr���d��9nY�N���S~�O΄&��5q��{��2�\w�����h2�k :��NK­��W#���A$�m}h�Q�bKX�&�z' n�M��-Ӟ\I\�'�a�ˆ�st�Yj#�' 3�^y��<y�m+��RQܰ�� q�\y���U�_��Q���+����>�Q	�'����W�BV^���^�`�ɿ��J p7�Ts�kT.{�������߰/�ck����������4l�f�ȼ4b�>W�e�g�Af![��~ѻ�0��{̅d���jr}Ƿ=Ɨ0UD[�<b�	MHu�<P�<޷��o풝���Y��St�j��WZ���>�3(��Y}^.1c��0��^�0��Z�o�����<k�uԶ�`Klq8�qw�{c)S�^�2�R�Bґ�t�HfPQ�)��ߔ�9���Iirɫ��K��ȹ�3XF9XXc��LՏ�X�Q5��d=n����H��Dx���?sZ�RTB�
��ѕ�l�ZOM��N��ӆ�o���9𫩢ǰ�˛��(aR�E�l[��k�Q��`���;!��8�U���F�ߩ�����@�w��m�e�_�n�V-�)W ߲��� `�o�ó�l��}}|�
�)c<�C_��-��_���/��~�7r=��n@�H���S��� �F���1^��)��,n���H�"�Sj����*+<�N�K)&#&�H�o.����`�TIz(�N�������U��7_��+��#���w���K���@o��$Rq�~z�.��#��ڨ-X���Y�{�2^�� ����*y�%
UG����D0�6k���FpT��hr:U�E��e�E�/�a��hzU�7�(6�8��J:�����7F�/y�ϳ-:f͖�<X-��-������iʄ�S�f?D���>���Ǧ-��v/�˚�D5��V�g�R�U�� ��^�n,A�f;A���������`t��c��i��&�2B�DQBd	�r�C���'Y�1�-t	���K�G3�W�H��ݭ���\h��D��W*���tb��&g���8��Du���#���yL��B�Y�������4MA�{��^Su����M]��^��f�}\W�.���?w���l7�y��W^ܕ���&�-��Y�����R�h��ϊ�RKJ(!e'Rk	:yl��c�!��*sS20)І����B�����[D&B��*yCe���qXu�<sZZ��@���돵�U���4�r�)�yK�e�ypl_Iw�%%��T�a��̫&m]#�a�~�I��1����9���;��������)�p{A���t��T�x�PLкo��A<�
�Z�݈
����|{��ݏ�_l�
z�&g,�~������iY���4��v��D\�c�oD�҈�cY�h�:�M�'_T��6��_� ��Ts��E�w1�˖)�rK��!w �F�C����ܡ@a��p�N��*~!l+ЬQ��J$� ��M������u.�m�9l>l�гY�*h��o�gfs�/�Y �\�o��/F42�r���Մ:w|>�%���.�P�^l/�[ٜ�|�lK�=��P  �>�o������Y�V �B ��CyxVe��sب���l��:/,`��K�nV,.}�����ߐ�93S_򻸠��%��m�z�Ho&�n�i'k��{��5��rY�5D�y����x�4`j�}i"�B��#���Av�[?��GN��Ͳ��I�u�+�NH�ovw��e�X�]-���כI�=X�h--��v�r�����Q��s>{���J�?{��h��<H��&�!מ��P>{=�k�L�h�&wLCnCmN�6��*y}�:�)j��լ}?�Vr9��Q�|�5�S���s-$c���8����j����m�4��-�k�H �+�<3.e������t��#5͇^V�/�{W�M�b�ݚ�l�c�T��tBr�u�yv�-�%��C`X��"$ ���LHi���:˶D|���4�Ep���^i(>�{����WRq/]��Z180�oqb{�A ��.��H�4��x6�f� ��VػSy	�wי~��u�A
Q�Ep����R��Um '�����.NkLh�c�k��~Sl�|���{o2œ�@b����=�N�6ڂ����0G�C=�,`L�msv<!��%����R�i��%�pL}}��'L)o	�Tԫ�v5п��8�F��{?k�\	����Bq��2�7��~+��gȧ�n��#������?�6B�13hd��ɶD��]���W[��;��*i��ڂ��	}�p�'���l��_0��2�5�N/��r�h��*�/�Y������y�Q�x<|f5m�wo�*�
R�
-���~�mKk����3D39�N+y���@����W�~�M����wߪ�΂x��7hs)+��&$�DH����ر5�7����3��M��J�y��2�7�'7�є�fg��n��ear�-����H��	BҹQC�LB�i��VW{Tu���I�n�������__LD��4V�i��.<&�M�����6p��c�����_�-���ÿ��1s��vV7��U�_���_�^�kNBk��1��\V'���#��8ق2��9t�X�� V���'��t��UT�aSO.�QA$W��ϧ�"k����&F�\��*v�1cN�/����,��Z��Lb "��o�:,��ǜY#?�˵O�Ԭ�$��0�c�l} ��C{c�5�Pe��0�H<�Qs���Jh?ښ\�^�Bӓ1�VKO�S����|+�N���w�Y���W�vk�-��&�M O���[gSD��(͟ԛ~>�:f!�AY؂u���k�J��T�5߆tĦMϢ2�vD~��Ԯ��&L����v���O'u��`2�rI��P	��-i'&]dL�Y��_����*�_1Hϗ�E(]W\�6�X�*�1���D�bϗ/9��vQgGIfDE<���e�[����;j�G�@��W�U��ߡ}�4�P���\4~=K���aW�y�>���ɢBxp��:�hP�X�5�.˗
�e�?����nS��N�=�~��d��B��c�Q'PH�M!�#�����2W�����B36��`�6J�}A�=
�Yamg�ݖ�Ѹ|Z}: �({N�P.��@��\��<%��OX�V�9�B�"��l��(LO���I�W�{8!���Z�:\����1F��k�q�R5�5�!�An�<�'�<|���=����P��/r^YDr�
�G�P�Bp�����Z������_T-dt5�W���������;�7b{@jD����'"a=ͧZQ|p�y[��͖=��c�]	3a����B`�_�R�l$��uZ �̚;\h(���q��I�>��G�\�Ӻ��jb���y�4I_���E".C�kU�~S��7u����5׫%R�mN$^2����9͛־<�H�^M���sz�+J@���ð<�P"�Gb����_ZI]h�ѭ�[�;�n)��~m4�$[�fa|W� }t+���Kc�1��O��d�sp'kv��G�o}��,��
�O�����E1���Rޜ�]��u���B�%X�Oč�ޚ�ȵ���ii[��5�(d���5�qo��� �r���_�M�����K
�	������5J�P��Y�i��5Ҫ ��p��r�laD�31�}�(Xx��I�y��A7n$`�h�6V�}��x����~�Hl/�Ҡ+��&|/��h�����ŵ�4����FU�/��护e`�[i6>*f�t���w�;}���D_��Xɳ�N��yĖ�E�| n��3���+��d��A:����fk$ӊ>��m-����¹����¨�BtRlϓ�Jb��վ�3ʀ7@�5��� ���$�K���@{��	�m������v�ƛN��+���$�;�߻�H�� �yۡ�+6S��QEA��APQ�wTBg$�8����,�m{�%���Lk Ҧ���q`*�Q���/U�kɇE"9kxb� �V>p����#��c&{u��Wn����#�����܆� �ϲ�d�6�D���vz��'�:
cW��0kХw����K�wO���͗����<��Ȋ�����i������Q���by+�Q@��~�!+�4�/���X��fPK~�DyX�m��wn/x�k�A��@Q&����t�_��|�dqZ]?. */�>F����v{6���t��`!h�d�:�2�������%J_��=$��������4���B��H:�=\e�L'���	���O��^���T7�k�3p+�҄W�6�j�n_�T�毫��d���CX�����/\p�Љ��w�Bj�;�)ia�D{��t��
��Ub{�-�z�(j>ȹ'4���#�*0ز{J�����F���t�S��s�C�c�FVQ����m�����`W���;��.��66�
%�x-�®_j�ґJ�����9��fb��|DY�!�:2j����0�z��pQ�Y��wC�LUZ�ak��hϬɶ�a�^Pȳ�SW�Ǎ��B��8�d��sO��:��$%I ,b�X�qʮfXo#O��+Ix��3{�l?�p$�t�kK�ڰo�0��]�V��}Qg"�?,N�#N��'��{�>�۰{�6ń�����i�k4);���Sl��&��a�VU_I�
&S�i��ʆ�*�5H��h_��T�D.�}�9G3/�{�)S�	��B������Ktc}����J�����|�q�g�S�O7�x\�)K���'j���1�ő��K�6��&"��8׸V�^t�"���!)��9-Ds�fmw�m��"C��ܳĶ��T�����铩�ta�b�9��8˙��Ȭt9�����f{M�
���ew��*llC�~H��t@UiS�Zk
�{�8[l癋�:��ďʷi���ٟ���7�Z�NL�=�;$��zd�dcp<65����[����V����f�)�,�b҄�*�҂}>��7�t��a4�hPH�[#�]���Q;��&Wh������[�3�aQ\�tj!�l���B?.��Vԇ����%GI�r���ڿ�8�A�y��_ܳ���j$n������Q��},��e8�صt�h����p�������$�Gf� E@:�4<k�ߚ��7�� �
��cң��v��Z���hH�_�# ej��	-�)��V߼H�d0(`]+o���*��X�a_g8X[��-.|۸s�� �P�V�$��{� �ac�hс}u �D?>��#	�%�/�� �p-�XA���]��='��m�0|�O�E2/*��00(3;�R��nWs�h��~  _h�J1a�B{-���d���~�Q���U�2>� �<͑k���;6lQ����X����
��)�'�~Fy�t	Ę����Z"����b���5 PWlkt��M�b}apg^��;"b'�{�/�&g� �Nx촎#��&�wbO�؉ޓ�p�r��%��2@�	���5�D�,M����v��H�0�qeU6/�$.�ߪ�3|����R�q?���ӥuix�kӲ�[�����o÷s��V���G"�Y)4աP3*�֩���T��,g�sxE��) 7s�a`�����q!=��c�e8Ir��=�_���T�QD\b�lv߽��X����I��ë�͛�2j��TT���l�]]?��������JY��pm+i��	���Vq��E�N�.�{�E������'!� >��4O�3�D@��A�������:ʉmw��z�J7}�.���b�������c���J��*YJD�P����z��C/K��/ɶC;���Y+� G>]<�Τ��T��+2���%(~jw�KS��z����O��|����IܕRB���S�8�^f��#̵%�/h�S4b	�iȯ���ӡ�!�R���M��d�D��ݶY5��{/�m@�b,�_�Rn9��#�e.���P����]��'���-絛]<y�wE���,HV��#��B�(�P��[`|�F<}��C�K��j��_<N���vím����Z%\�|��|���՘X$�*�,���{�B��{P'�a�/�*�B�C��̞���EN5�f�^�DW�:@�2������'�O��/�PA�%�P�aKW��Ku���~�&]l	T��� ��{Qٝj���B�,h�&v�'ٗ�������٧��4Cm7���+)r��<��I����0|qֿ��:���}�S5��Ɣ����<�UoE��xWGo��z$_ս�Y�ԉ���)�r!�6P����$���I0z��� �}rf9�v3�1/x
�:�۳�C鶣��ɍ���h��sy�O�"�[�45��8Eΐ���#�0��
�A�^+�%�w��Y(]Q�:�x<��K b�[�6UMW��^��my�ʸ�1��m3h��{�)��}
�b�|���:�Y�ʰ����G�0����jg�`�x�v$��d��{�����]�m�bc:�s��X����(��R�Z�����*�1���i\̋˱�f~ʳ��Z�	��*H� ��"��_Z����*�',�z-�	��M�c^=7��V�ǁ��=��� �� E�n׷O�[�^��ҫ�I�������_,p�n�0���sS������2�b�N
�y���`�cֺF���ʌU�, ���} ��*�1(��-�MU�|���`au��ԡ��O!Jm:��)�C���o��u�H��Rg�1��X�N�Z!�ܸO����6�t`�E��b��^���X��
����?����U�@�D��o��n�;bN鏮	Te^�Oix1Q`b��;n�=��h:���9䚓���żI蓌��0��p�*]�t��LА�@+	M!�AHB���a��O��c�0�A�����UEP}��b)��0@3\��/�Ez�(9���7���I5	7K�{ķEv0���0q��1��S.X3�iWxj���H\�8�B�bH��N���w�]yٕ�r��ƌ�l\@y����G���KF�*�9J��v}_��(us����E	��6QC���l��|3!�P/ڮ��Rx�F@��s��`W���ى+���W�E�8��-���̃��vH��Ạ�޾��g�J?X>���[��������v���wLQ����+�۪lY$��!��X��c[w�1���|g�;���UQ���?0�F��<?S��w{0h�<w�}[Q7f�bպ�9Uѯ���H�d]�Ύ���[$�IK8�Xm��/$l��N�t&� �j�i6M��E�EcahD�bro�b�9��,Q|��ݰ^���n�Y@WG�v�u������]dmv�fNT�a<�������22��J���z�jf
�%����q����\A3�p��Ԙ5kB?��	�y��Vu2���H'��X��_�d(��<�s��s��z#�Q�8��EX mnG,1�z�hk�nU��(E߽&DSC5+8����#��W3r�u�����tcrU\���̥�uj�dQBޭ�c�k�q�X�8ͯ�á'��=l�r��t���^�������Ȉ��S5xs�^ٗ(�Κ|��ܐϠW�>�}.'4 ��N4UY3\�2��<L�?bU��&�"���4���~a�s�w^��$�^ܤ��3k����[����9P��L�t��c'���;�m��c��Bu��
��.��%��RⱀJzx�5�x��}P����ɚ;�Q5</�Y���A���l�I��䋗�DW=�\i�p64d`�~C� �W��)�0�j���=��L�bG�',x53�V�e�M������l[�na������ӛ��b$>ɴJ�L�.N:}Ќ��W�҉�"�{`�0ΓȂ+�(gH	�9'Ž�=~�	p�#��A`�5őj�d[�ʹ�p���@����
��eݿ��WBCf�oι�Fjd
��b��r���>�aE$G:�lzݪ�<�.�iP���@��h��R;�(�H	��a�K8ߺ�OF�lߖ��}A�X��h�@����"l]���3�Ӯ,%��� c�>������2���g�Ϭ��ϑd2�������EC�=���-ʢ��=��e����Ҩ������BP�栃���lX`���k�q�� %��s�~?H0��kN�$�&�70rf/�g b�2�]��q���D�W��� ��C۹�]�>��ٯ�o�h��k��|~cT��e^�~�-��4�^M�W�0�~<8��p��^���6i(�R�Mt�H��t��u\�CЧ1�2�&@�G�~ܹ-��ׁ�qz��B5.�����n8^�|�d�&�۟�Q�yϦ ��2̢��jBx��y�� ���F,-m����tl�����%��I�b��D��rC>��ղ��C����]�~�{��g����<�\m��?{��4��X��.�|�;"q*�7�Pb�	����=F��N�7(��?�έPW���1�+vC
�<�P�,߾{o���[d}n����V����W�>Jk<�	;��b��K�z�@D��\l7'�$˺���4���M薞�s��X����Ck�yl��r�^lJ��'��DV`�'�8�g���x
�������7��+y�I�h��`~�o�n}$e�t{?�z:�
?a)�UNDs�V��ڛɍ�QR�A6���%��O��,�p�$,v�%��T����%,f�dL"Xs�*7/�����T8�"�w�D��̘}u�B�Wmru�}�^�v�s�2����T���SNT!vZwL��v'y4�|SQ�c��c�c�v̌�a��T�%8Zp�M�4�LZ�cd��u ��nV$zP,:�RJ�\Ӱ&��<c�u��'�Ip@�x	��9&��p��i_�T�8<�j8�ͬ�-� ��L�3.�'�l�f9�����t�����4�,/�T�i4��'e��L������ h��R�ܽL�xV%�T�f�t�����ԓ�f�_��\ ��T�4�Z����#�T�I6�����{������)1;X��e�()��>����Z��&�`��y�Y�/;x�?w��C���]O����a�0�3Õ�1ذt�6v�7O~߲c/+�5��V:W��K�����ؼHr}#����	\6x�%U]w�o,\T�B��,�"����Za���XT�Z	\��@H����2��y\��(_۲Oq���|��Op�<}}��/����"�lĮ���a8�"#��N��Uyo��>@։�ۧ�#}b�j�=3�xg��BAH���r}C�����s��Q�BT�p&�I����ݣ G�G���>�0�ב��gR=���uyKw��y�y�`)B6��͹�`y�JB�dJ��y��h���}2�	\T�J�КKH�OO���Ş��e��y"+��J݄��]ثHݫ}�<�P� m��l�|͍�a~ۿ����x�𨐴�ˇ�Q�8���2�]乷��C�����;$����"��Oyr#����ޱȅ~��.ev�o��=��i���6��l���t<&I#�\��(4�yHGP֔z�,e�{�WE-Ɯ�����z%�X,'�U�fUt�(�A���>�à���Yu(�)C�4W?GЮ��mN�Z@Y���3��e�Q���\�T_�JI�ψ�s��ҥ1-r6���g��E_DSܢ�����J)"�|N���z �&aJy\(�XWZ({^�l�.�j��4g�ƥ� �w5�O3)�\O8�DC��z�b��C\����ҜQuq���p�u��@�%�T5�h�Y5++ݡ���E�'>��7�D{��1I�'#e���S���>�E�5Ҁ�0�(�;��fש��PN��׵bE5��D�w�uƹ�naA��"Ӑ�ǣ�of^�y��P?t���u�Mu����e!�G�QU�M�][��u7��ѻ�k��"��ʔ.P�%�UȊ�<<&��
xA��@E>���Ob��G7^�(C���ab��@��C׏���r^6���R��!5�U�A��Ѳ<R�ce���L � g%j
�Ù�t�:�ȫ[�Qɚܓ�d��|Qd�@tS��2k��Տ�=~v�y�C�j2e�|W���V�^/�@�&Þ9�d {�7���M"�N%SHT�q CS�h	U�a���s�h�zവ䩁�'��(Sy��48��j~����b2	��,��鎼 -Y��r?��Wò�YoD�	�+-z$�I���{2K�e��ΐK8Ƿ��p�<>�k�}�^�*8�(�S� ���u�[?z��W���(��Dz�4�/�G����?��:G���1U~���_�cTN����Фcjsd�d��Q/�cS _�'����ۿ+^����݃"a������Z콾�E_����Y�z�)�c��Ȏ����zQ��b�Z��Y�!�GV��+�^�!��~��SX3���,ОfǤ�e�z��'��.*�S����YQ�6��b?wy���iP�%t��u� ��9=���� ��o{9Zd	�R5.���s[L�R�s9��߄��w�/�@�I_滁����V>�vt��H��R�c���PV,�����p����з�ܵ�/��wΐAkTnT��	@��_�-�y��4�lM9�2�z�@y=;�#I�?�=��'?g'��쵲�^���M9@߰܎u@Lz�����y�u��5k�&�2(yKXEO�2�2�)fx��H��t�3CE@��z���LG;�P�A�Z���b�������܌��T�Ş�)�?i!'�����3��53���]2�7���W�V\s��mZ�]|�-��}��^c�-�t
��]����K�
4��D6�lS�DN�,�y15�p�h��PW���vL��	��5F�VS�X�����u1�+"�gÍ��A�X ��|6����܈��T�t�F-/n�VGS�Xʅ����&�Э����R���^ŀp��YؘϷ�u(L1A�f��O�n��\�u[�K����xB\Ys��b��}|i�v�R�=)�%C���n���g�@ �v�|C!e���q*�m���u�xNT�p�|Ml�Pl6��y�H���]��D���ID3^�+����w;�og�����HVJC�t�Ed f\+
�/� ˧e�5�J2����_rn���悙�'��`�4�:�Gk��ԜWIK��r.nv�H����@��Ɖ�2��������"�L����?��%B�gB��Ka\0Ē������y�aL�<ȗ�=���n�v�>H���AMN93���#�o��}r���£�1���)�fV����%��ƺs<C�|ۊ�>�=]I��?}�Y�_���ʺwo�Fջm����dr*L:��K����p�*$U��Xv,u�xB�]y��a�B�����e�-!�g��.����nt��Z��kQ$@�uP��il&�3h+��$\�x4t������\�d���R�?kY�Y�Ya���t�5��)_�;�hgS�O@��a�2*s��9RF^�ͥ��w<u֡zx�YD[SNX4����#Ug��v���>|�������#:�V�!b���3%
1ٯ��wVK�Jʚv�����g���h�D&� g ��T'��c	�[�	����߅��5�_^nϷ�D�h�Þ��بQlv� �ѷ��|�Ë���74�V�.�hZ�0~�xC��c�1�k�����7����=�E,�s�R�oAloSa��=��'�$,��p�(��X\��������_0����c�C[7�%V�&b�Cf�(?�r�Е�H,�s�o���j�����O`L�����^��hȴ����/@!�����nwo�W�?UJ�q��!|n�=vo=zd헌���1kH�\�kj���O����S��[�LL1}��[	��7����<��-ʶ�C]x�n@�E��l^�Z�x�Y��-��b�`�U��`,D�^�թR=Qt�SC�?u�|[+��Ҟȫdo>�9�ߌv�F@9G~IL����=,'e�k��w A�ioו2 �xը {:�*m%p��|{���B+�B���C^aoɡD5���f�5�#�@h'���1����e�ԉ�*nr�G�*7��I��g���m��8%�������I\ms0����]����!E�C�e{��.$��E~���sd��$�\��z|��3�ɷA��i�(;q��E����1�<�IvИ��k�B�y����_1�#���R���0 )����@��Z�7�9M�� ��須0�4Z^�!7��%%�+(�!�Z����ب,^���������H��Ky|+��Q��zx�3��\��9���'0r�ƾ�@��1P.!B�>]�2��P�Xv�Ⱥ����j�Zf;����ړs���W<�F8�\�����s�A�����PoE�Vs`<�Y�{��*y��	����[1�uH��u��GWg*���|��֘c�kT+z`����`(#�y��2�N:��=��x�[�\§!?�l��[w���6����/��Dz��z=E�Ż	
�!f�6��������:# ���S)�����_C١�4�5�P��U׵rE >���+�fN#)���XB2nFZ��P߼�]�B�X�� � �9D��T��aY[bw���[SI��O�V�X+0�g�h⚯����.���� ���h��mrꏷ��$#�&>-K����_#+=ԒA-��C{��7	�z�;ȁWD�~��
D�C�g�<�^��[��KQ|$@*w��B��*o,������E�BwPe2sS�hE����4�$��\�]�%�+c����/�W��RZ����-�@X+�F�����s�W�2S~:����٭��OO��ؚ�\��>�#<ʯ;��vZ�����J,З��H�ޗ���!�>D� �!�v�;�D�G�Vវ�hj6�h�1ɢ"�bC �X�E��C�V�� S�E���v�|���|x!!�+�ղ�]���ATf���s��,��)�V��!����1���&i �ܼh8��U��J��o�\�_�(�W��%<ם��O��;{���F��݂W�S/g0;�zg�Y����0��-���x#�2�����L1d#l Ѯ�b��0.)K> °����k�1�=�4�3��+a3�f~��I�3/t��М�🙸�s�	�r5e3vĪ��e��t1
�~��c^�TU~���ܴ��k@�Z`���ם�)�������(�(�y��{��0��ySt��~��ps�ظc�SA֚��?�VVݰBq�#��Ҷ܁� �e�>�)o�:�_
b�kg�9gl����R�I�a�;>��,��v�]���@�YR��v|H����2?�^S��}~����7��0�hШ�,8����?���fcV�P�8ݍ�	�br;o/�=�ъ,�����ǝ�c�g��{��P�s ޹����(̜�;�zg�{P+'�N���xu	c�h��F��Oc3���^�����qo ��J^Ԭ�kL���ފ�%A�yIq���h*B�����<�ˮ�p���'a}1��M<	

]ޑ�����j;8W�/��ux������qπxt�C�a/KxhK�DZ��u|�ŧ�xyi�e^5���ˀ��p_y�O�lalW�y�n��Ok�]K��!Y��BK���H#j��HPGô2��wk������ɮ3x���M��v��@�yL8˔C�<�F�K�
6Ԓ��D������m���m���OS���Q��|����0�E��f5ѵj���
����j�o��^"�x��(�O9� ��Ь	��?^z�������g�<)	O՘��b?��h:�W��ï͚�)r�?l���cܠ�S�P(CL����+rLӅ�8���.���g�=P2T�$u_������oq�hH-���Y��3�V��UK�ҟ�v<Q�-By�C'kY�9k#��#j[S�|髥�~�e��.���K�l��91	� i�!Z.L��>�_Ύ*004Y��
���6��t2��db��h��Ӊ����o�ܡ�q�Q
�s�C>x�~J_�d�=���Qm��8�B���jC��k�x2�=u|��\R�g�!��L��U�h��l���$�����[��/�E�A�, �����-3i!Լ���L�cV񏤽���m�� �������hj�|X"}�uf�O'�3�td���T|a\��\FR�E��Y�3�'Z���A����,q>�2��R�+sE����>�[K�m4��Lh�Ixz��{�j���E6�Hw4�}n^��:�(�S��v��a|<&)�%��R�D����h�DtZ���` �θ'���wƔ%M�v@��U�?a�>e��B�
��K�F��BG��"+�CR%C��%�l`C�P�m!��m',H�����\��7��}���Feؒ:"8�4��bTO=V1��d���y���K��Q�h����6���wR[�����:�L��m�^_b����<|,C��ɡm���!�l{���U|�#���_M������Qc��U�A����َKM��?�A�H�.~�6�t}�/��@N�Pj]Bm�D�����WCjk���#��m23��!�E(j�: �������r�"�ډ	�'�{�4�9K<>.8���òd�~�O3F�A"���!q�]/T<��8E�W���!kE�<��V_\I��c2,����PѤ�]Ʒ��L��#D
�/5�%�L�|�L�[1��|��~�ڱ��Z0<��ژ���F�;�`�
�4s�Fv�����Ҭdȭ����p�CR�X��\1W�n# ���TD�n���:XТW)&p�b�9�Y����	cR Ք5�_J��'��K�!\�$V��*(�ȃ��L����b�0&�eiE�f����'�f2����iQP:��S>ʝ�]�Q%�wŏ�R/�5�+�v��:p�u��R�!�M�P�Œ���+&��>ū��{�UЂ�Q�3>㼘�c�[�8�"�Z��('����g��#q��c+y����vU��h�^��ZHD��(\H��Մk@��N��<��~�mO,��%v�s��a)O#�(�x\�I���8��,���`�D5�L����sv�U�Nyx�~�X��&����0l�ou�\s�3"��<xW�x�j����7NH�&�!=��n�[��� �!��}}�2�ӍQ�3(�xo�d8����$A���~���I-]ڮcP$��2��#�_塾�q���?`b��o�YӠ�T�J4�$p���Q��w�����XAQ Ջd��S����I�6��+�bf�>h'�;����쾰�@i�X5�._�8Uwh�)�a2I�0Ι��.rh]�
��%դl�p{C$i�:g|��(�ڹ����[X��
y�Mma&L���l�z�j���fC��n^,zI�l%{Ѷ��ڏ%��NAA��;ʈE�Bf���_sܻ��߃��Hf��g;/��-g�:�w�_��"T��p��Х��t��+��	�E�`c~�w^E2�|ZQm�Vak�+�L��䶓�AI?u�P�aS�iu�ԫsyD9'�"B��1?��_��u!�B Ao��D��x�o�G�Gِ��[�ԽחR����d���<ipl1�#&EV/�I&��k2@,�o����w��j��ir�|�+܅��� �rX2J����va�k� �&�'q�i̢_8F	X�Z}G>6�	��m�1ޓ����oYǩh)��|�b��M�Ğ6aA��"��:��=E�[��團�+��S<� 'a��5�R�6��H���y���vj��]�Rd�f�!��X��0\�%�k�\�*�)9�(Kq�Yve��C����Ğ���{ʃ^��>�b��3��;���ɻF�\�D�*X�F��I��>��U',�p��_��pjٲ
�����VF���2x�H#���@�jU���B�Y�ޔ��5,9�Mc�Z���4z�.c��f��{\I�jUЫ*X��wG����9�������gw\IU��q�{r�U�W�fn|+a�f��Aͳ�IY�x��`�܍x%�R��l�׷M����F�(˸��d�UER��ƺ�|�X�It�OٖH�Zy`��hƠ��29�B��m���~٦����W�T�ur�W�z��� �
�([� O+!�H$ �x�)�[�<�@��������i|�$c(�#�����P#����n�&�+��<OD.����ZʰkN�qy���������7�a��z{���8:]+�^	d��(%���B�t^�|���H)���Q���9H�X9[7��k��`W�猬��*�ظ���V��T���/6X��'�G prYtwI���2Z�vos�J��}�`s��2��1� N��Y���\3����@G^���X�+�c�QW ������SQ�M���!ȧt�I�:��Z�{�h��\�S�_D����Iw�t1kc6����SV̈́�Zǚ�F�Hc�E�l/n[�������0����Hm�?0���>�Q֫���{aF6G�l��PȢ~XHqrΚ�\2Mw�R�"[�qm��/������a�9U�_sr�� ��R^/�'���*7�\i��ę(��T#�
ِ#	 M���ş�%�*מ���\� �[7�"�"]�}Q=eyw$0y|�b���	p{����~�+��TΕ�ko>�
�%N3̵3�7c�7m[�sN�dK�3��L����PM�U����yK����Q��Ԃ�q�d4�j�?���U}bp��w�%��@�K�[wN���}�FR%���K���4�����˔�R��B騍U�x7����n[t�#3O��jQj�J�S����y�����b��	� ���	)	?�%���@�Q�z����N��PH8(J]U��i��Pj����ӭ�j���eŭ�kN��{�o����9I}���z��Ҷ�@��ʷ>�ǈ����e��U����Y�"E �g?��Ҕ���m����m�f���1�v�|͖��B,�`y�M��wA�`i)��{��w.6��D�̓�u�ѿUb�;+�E���P�!���H�՜�GY��]����c�׈�)�TE|�T�AGl���h*�'{���Bz����f$���M`1�`��p򟍸G��ȷR�i�^�F.nc��Q�ZJ�`a;ITN��Q�XOo�F��g=���ԝ�t�����2Lz8��m*yF��ƍ���A��Bi�\�4�?�+���Z���N��!�THVspy���GVyR���[%�a��Q��TЕW�V�l}6�aWk;��2�7�o�O��8�m��+ޢZ����X��*Ui��|�XlV$JHV\���"`!���H�����t�� ﻁ<ؒ��P����Vt�	V��A�7�a�ꎸ�i</�ʬ�HGh�5�^��Y8��=���'9�8J}��G�H�),GE� �ɹi��>�j,�T��rAϼf��F��v��	?2�7��J�q`��ő@�D1�-P_�K���O0ި�d��3-&���U=[^pe�#ce/b4�9��q��'�to�PX~�Kd\�G�"��`RKhQl�	bAn�{����&�TN�T�=��_�Ђ�!���to �*��.�6�mܙY�p�>�A��0��od5i/�Ҁ����,���7���0P�p��6�Q�JQ���k����/ZĨ�k���,t���Y=� ps�4L���=VǄ�!E�����Q߭[�&Q҃XЍFN��aO ~�}.�{ib���G�;)��� p%�w]���:�pɎ����8I7����؄��q���ꤹ�
ү�=��A�0�"����"��i�9҇�fw����7����Э�ё�q��FJ�,�u�1J����8���_fAY��96�`G��m ��X�B�Y����[&t{�*�}�9�ܩžb����q0���<�  !�)�4��5�� �*u@�ò��po��/5��L�}F.c�B���� �g"%��L#@��0=�x����e���(V���aSC"r����`���g ��{����O��y�F�pk#����H�LQ��z$w���m�2]����J��=��W#+�۫Wd�[�. 8
ԪH�ٗ��6���]i+�����I)g|��'`����!��*ZW�����c<4���+T�a¾�m`�Jڻ�CyW�,��8�0�r�>HU˿8bXQ�Uɒ�-׾u|޷Ao��{e�0�o�~�P��6_��'�k�Z��e�G�'�K��>�J	2�jZ�qv_�9���]��N�G(*ף��׳�W��V�����˱^���m��y�i��ڝ�ͣ·��Ϗ� �t�nn�O_	��$�����t-� �p�%�l֟�7���LS��E�jt�~`��\z�ju@�6��}w 0�F�OjS���CY���m��d<Z�G���>k� �k�t?�?�)�:c��ە����FP_۠~F�B��_��4�{y_���Eq˛T
3��7y�/	�V�h�!m�ʔ$P�Y�*~z��T�@�V�L��
I�*1�e,:3����I��-���;���}�m�ߝ˒3k�ғ����6�Z�G�{X{K��/�m��C��b
Y�Ԓ*?��U�>�U�/{:��TRi�p.0�0��J_[�9�d�͝}��L��VՉ�r���(����?��!o�#U��S>�jv{TC���,���O��ۨ��q����ڳ�<���D����ۮ���h�@�I����E%ң޿a	�����k��nz�Si��h��p���{��7o�F�Jb2!�BY�q��[��d#�j-��m?��=�Ņ
{�'$���i�%LxA����D�&M��9���9٧�B������4��2��Tӕ��e�#g$�[�6)/X9<u�H�N�o�q���F揓�jj%z$R�	����~�����2Ej��_�e����*�j�-�� �Wx��V�L6�,�z	.���_*���BZ�pi�n`�J�:���AW��L@��Wj��w�M/&��PW��`�]wyFf�z6M�G#cmm�E.����+bLqe� �2r��J�W�k;½@"���gwvZ��C�:��2���*\�L��c�	#�E�}��Q'ht�Z2??�{_�������>��,x��+v�o�/��.��nf����e�@_C��^)�$�J�\s�l����W���ܱM|Dy�Fu�'�8��˘�2bi�_|j�;���6�m�h�����F
"B�-E*&�
o0&�����P�9΃̯(����@�˺�A}�a`g��{�	�k�"B����vUȵ�_��c�R���(��X���	)Ǥ-��XJ�;�Y�鞲ڪ�[�̩��.�ςIT9L�yL2\ ���Y'�F�>ň_��Fc� ����hX	�D+60� (P}uAV�r��wYҔ��	�]]Ē���j�Fi\$�r~���p�n��s���9��|��w:�r'*�"ٳ����Н��N�Mx�d&�\�Jv>P�3�Oة�+#N���m����W2o�'�rO��E�T@�W_3>��Lf>�6�1�J�$E��AD������i$��'�Ci��#1;�Ҏsr1��=j���8]+"��ɖ6���� ��ԝ<Ad2@����<A;�?�����w0>�)~���?��`MN�߼7�PS�R�n��d�z �W���a�N�N�ʡ{ۤ^����^j�W�E�t��"CH�HU�o��o��2��e�^J�r�Sec�n�Lʼ<M͸[6T�;������I�y�Hj#u1�##��B�G�!��nT���5�p�W��c��� ��d�� ��
�o��/>�pRp����yC�&��| �N�U�
��(� a�Cn�	�3ؕG��[�a���۰��yC���Db�4��5��?:��ǖ?o�1�^'%<2�z�^�蛂����EU��E�z��NnN�1{� ���	��-f��"�˸��kO;dʘ�QY>�)3hj5ns���j�{���Z��;s=g߲�eN ţ�km��Y8���(|7E�Cp�Nj��b��_}k
����D#���[W6@��e�
��h�v9�pg�-�	�l��^�@�������-�#�
a�Mqa��(��Ҵ�F9 �3�����x��ط�D�>�R&���T�y��v!��$5����7���)/�W���y��Ŏ۱g�����`u˶ژ���r��Y����Z+�W�����$�;9�yʒ泥V��V9�
���� �����ʪ*�T�y1���~
�j�j	P��+���i�,�F��T��?lU~E_�{��燤�\�i��y ��#2ch|Xy�5~q{ƺ�d��0�&09�d�c?�}c���m1����p�b�^�=�C8��!ȶgmB��i����a	X��iU�~eP��:1�u���$]�?w���%}#����P���Q(��L;�َ"�RF+������ּb#`���o���>�<���W{�O�����|�`�w{.�ΰTPx���<Y4�� ����M0�!u�N��n�c$�:y�A��^SR��G���hI�/=v��W�W����$	G� �Op�_�β�0�ej@�)�b��,�5�}D(���Y=����u0�|V�g��y�>I�];N��8�~s��/��0�Y���q�@���?���Q�w"ᤕs曁f#��.��f��m��斣�V��+�ҪI���߷Xs����t�:�h�KU�EP�lC;n|�Ũ.clQ[�#<�B���fǠ�o\0*οVm������b�뉆S� �9�1Y�'�m�d�/!a�a�NUr3\��O^���մw«A΢]9�ෝyh�왦L�k$���/�vn����xl6_Z�҉�ь����z�`2r��H;_^��G���~k�pZ�a[: kp�b�p�D��
��S;�MFJ�o6p O>�F�t��6S�U��cʦ�-�Rŉ�D{"���6�&���� �<����/4̼gF��U�`�~ۑ�ר���_)�i��/�Ի�t�S�$�z��|�Q(@��ku��M)��*���8�T��9_ց�K��{��H��ъÜEl p]����P9�]������"�~���aFm$��a�^��Kg��NYqA:�@j����U����G��������ƃ��~��++�H�G�/
�H�������-��ª��*y ]����o�5��a�!�8T����0qOx��/%�0�B{��v�b_�I���K%U����tl9!�a���e�mp= �V���W����F|�F�.�^��&�;m�C�a,]���;R����?x��c���K�6_�����0c��׮C�)w��r��?ʕ֖Q��Ʌȵ�N�WhIG��l�����-�d+w�n�kA�1`�{�2�6��$�A�v��=��a�1����M����[:��&@�թ���h5C�dY���0;WSB�9$�R����9U�^E����a�8t�V<��]��i�>13��ʾu�)G9k#�;Vb�� ���L?~�Б�D����kGj<��mb��Dd k+�bcI<i���(<<ɓ��� ��.���
ɶ�
���!]	#K��f(�)R@�Ö�DXi¦�0����>��j'���/��P8HxU��N�$��QN�{-��3�
�U�`F����HW�����=�;�&��:�$R
ЏRϥ�@�s��
jY���tx�=�#�(1���~����n�@f��rK�� Ox�� �X�;��1mp7�N�n%��Y+�Ѭ_\ fx$)�Jy-��-hӧX��2�~�+[��,�Mo���'�RO�â��5� ����n톨zqv�R���~j �g��ŀͷ]n��LtM��3��f�9�3�'��=fm
��>���L����7�P�����g!�3�^&y�[!�s���J�:t1�����\�p��9�Ϝi��7<�M�0-���t���������`c�1�����v�H��%���/����!n�	Q�}73r�o�H�K���a����l�w�K�F���P���b.�O�m`o!ti���Bf��߶��[�?a��pP?��Gu�qؔ��=�&q�P�Ly���4�~|�5S~&MJ�藍�L�!��֜�ũ��(K�(��Pɬw���Q��dz��dQZ ���^	�i�
�/��u�)��XL��z��	/�.>����rK=j'u�Hfi�杣#�a�Ł0�Y����m��IR̦p�ϵ&��_��I��n�3���}"a��m�P�,�K'&6SH�z�Z���$=������[���;��RX���0���/��/L=^V7�����j�����;�����u��Ʀ/��1��%F���%��OC�ߣ�U��uk-�TT��a�zx��H��+�,Vj*���knU3[��\��- ����-�L��&X���3��c������Z�8��/K�����X
.T%Z�{L�U��y��l�Y�j���%\���`h,�i���RLͳno���﵀��i�����vB���ǫ�~�|D|� +���0={�Z��@?��D�pH�Sɬ�(��p�g$�+�M=H�5tNFߊ��У�,�\�@U������-��؁m��|¦�,ш~��qh����!/�ȶ�4�����W͜hY������V���'�����y��_���	m����)�^��֠�N2����> 	˂H�ػ��(������^J�a��!z ���邶ѷ�ibYj�U�(V��?��HS!���"n>s���s���fW�J?w�E�3��3�Q�� 8�$��Ƥ	���b!i&[� �pk]Q��r�u�b�8���:�"�5�RI\c���P�E�J&���î!��t��ħ/I.��k�ɥE�,p8�X���Vq+ǉIK���/��{p�J�P}Tڈ5K�m��R}Tn,8c=F0���=K��5R�����@M�f�"y�+ɹ:)z�~���T<T���$AK1-�nl�j?���rM(8QW��C�B��\{�yR�W�I:�d�'�V^��t���2��R����ʣ6M�D�oPNW�l߀�ӗا��a���k%����L`N��D ��	�t��9«x@@����,�V'����`E��l����R.!���{k�n�ߟ��#N�6�u��z�s"YE����u�#M�o�E#_���ER71��m���N��?�������b�������������5��},����-�€t��|]�����ٜ1F�3�I���&w��¤�nsQ�����#��l�;�>ݧ� �{���jߎ��O0c���#��;2�K<�Ht���2��6K��7�,��a�<8�">��0a"n_b��@�ZQ�o��8�x��1�P���CB�7ϸ�N_zZ��qA\Y�v����8e�5��͒�j=!Cc7.z�5�'���נk)�O�ջ$j�Z��p0����z]k��y�<]U�}N>����+����I�S�%�h+ �"3ʩ�]��z$)�`/b�(�h��$��S�C�r[!� �V�0�)��*��	a� ,��a�*A��G:��/Ď,��`Wɬ\Pt`$N�g�KH��U��.�<��g;�xa�mB��0c�8l��N��A16���=jEF�'QN�����)��x��E�A�sG�֍�J�u�t�&W���[k��)7�)E�}$,��g��g�j����I�U�6�8���E8�Wޛr��e6��t�E�KY�L���|pM�^.�g�6�ܙ��Xځzݎ>����i��פ��B	�p`xT���)�E��$�*Os
��9���O�/B���L 7 ɽ��1�j3.[\���� �"���΄�0��3�
B{�"�k��+�����crhk�I�Xw�>C������+��Ý�ց��L��U�.������]�]��k?M?Mty� �3�R&�*⒊����8t�&.�@^��F�}UGA"Y˘��n�l�D�	���ml�;�B�EA�'�E�-N1A��O#ǳk�2��H]ΰ/�t�=3��)���ix�u��O����ΔW�V�����X�R�� F��VU$�Cj�.�7o-��&��wU���$a�\�c8_s}��j8	ܦ"M�R�'I�?|e���,^]i�-�w� f��N��m	<:�L�����9xn�l���C`�FzB8����Hcw6��R��f�D���O�ok��n���Ӯ�O3����&���2������~b��E��%K�������C�G�hy�iQU�i?�J(*V(���I�6\ʐ�mb��&_B?�1����2R�
L L��Ega=�<q�y��揭�]��F�-�>[$)-�<�%��
�>�qf�������cpi�dD�y�e�a������n����.H7�´��fS�Q[UJ���Bsꍮ
v�� �QG�zEV��SN�����P�	~���\���OxAg�U=>[��.���o%���Q�'�USb�ς��M��	�HH��+��QSu���|%7��g@�-+o��c���I(�[����r�٣�u��C��9��$�2��� ��8��>M;©���������7Εj��r�zA�#��U7�ą�qE�6Yôn���lܻX���[N��z���^*�FQ��>����8�{~P�{�D��?`(;g�4��y��Kk����:�R�f7l��Xt�7/R �E+�ZnCK�1�O�_𦗯:���i�U���Pg�`���:��U���i\mH���b�ʹ`u�3	]rq;�:
�N	���2θ�s�{�Փ=���5�
���>�{�1ʳ v}{�;�-j}�[j�~�	������d����>=��b��Ͳ�!Qf:1F��eu���̬�g�C9�p�M�[��4�� 	·9T(,�������������v�W}�<�|�ŭ��#u��O�9�ұ�QC#�m�k!����G+%�N˫h�j�k��D&��~@��%7���,J�'g����F6��X!EjAHx홂GI��sdf�k�O��VN�-��z�q��� �P%u����P5��ɋB[�U��[�ɼ<eش�f��Ð"&"׌�7t"��������<-%q�(zb�$B���$0�����-��t�o=�zG���vY<2��\�6V���,L�uJe��+B$!'��hO γ4Tl���v]t+=���ͥ�
9�9���"�Yb�ɗ�W�$�.��u�PMZtcu�\bD�	7Zsj�;g9,�Mأ�� hH)~�s�I����#�(����
}�_@�:��os���05#��J&��8�-Y-�A1d�i�JsG5e��^z�T�����b��jS�8b��Ҍ�1Eǵ�K.g���CI���]�u���"��!�t&�I}����w{�UeR��@�2H�_���m5߹zݰ�{��D`Tm����DB��"�sJ�f��L:�\�)w�m-/�QN����o����~���bq�]�T7!v��j���%<o{�ۑ�։�S��]H��}ɬ�_yp���a�.��<�������ѯ����G����k��P'u�cs�a�,��ݡ�ޭ�a���r�(eDQ:�(z������0�����N���܉��uJc���ǉ���>�U����[�#�ꦈ~/^����"�5�Ylx�>E��6���Zv�,l�u,�ۻ2�Mӌ�r#�F��6I�1� ��o�)��Z)�CP���	Z���Ȉ9�3�I�萊�Թz�3�A�T�wG�v1��5��.c}|�?g���g�4C먲Wr�5Ϭ�U��n���"�U��Ă�E+Yq���R�ڼ����H�?Y�>�����!�K�Њv[��U�Or}�Je��-pDo��ۼP��&�Q�Y������s�z����'7�Rd���Z>�4Ȯ�7�n<�j��]19��G�(�U':;ހ����*�&����&%YMW�G^��2Y_ֹr�?*�&�:��t_������S����3JB6��Ļ��|�����2�J"�-ǔ��0Q*�ވF����:�:[H���׻����Hj�LH*v�PkI��_����6�	�o���׵{� ��s��_�M�V-c�B㏍̃<$�!��_����z�̺L�*��F<]� L���E��Oe�D��jU�S^�A>�^ï�	����~��T��Y�=+���x��ӎ3WuD�sT7 �ȹq�ͱ�Z����J�����U��l5g}��I�p�'A�Qp�����8|�S����_�U���/�5 ٰ8����^�����] 6�^�J����:�¶	g�/�գh�[�sEK(���v�d0���+[J�դ������M���5v�-|�mp$fA�=u(��r�C�Ԓ�«���~t�ǂ�*К�u>��1��p�>������:���	�zhNW�s����0��٘�v���®X���Xv��#���s}N��ʻ�V�����b�HT!��T]�/���[�h������b�E���vG��&��f�?6����G�_�痘�zYݐ:ax�*�|��l�V8�e�1�E����_\���)�ާ�	�\y��_۽L�R|�����B9ٓ�L����Ui�Ӝw��/�����/~S��_�
T������-�O�m�� ���ĕ�Ҝ\�����y���k�I�y6Q�/�It���m��y/�01����J�}�������,O�J�ᡟ��Ӂ�ྲs�ւ��S^qЎ��+ԯ"C#k���c�?xbp~�����qv?z�"1�K;���b,Fñtj��|�	Ypf̀y�]��h��p������ZO����k���0Os��ɋ�d�m�;Y�B(������'jm�0�f�(��:F�F�D,����^'�����u���G&8�]xy��ݖ4#�i���1�1����</͌;N:-���GԾ���'��ߌ�~2�*�u�e*��$�n�F�弚 �6+�^OM�/�����Zjd)5_]�u�� Z#eY+Qj���jj�AL���#����X߬�C�Oo���A&���m�}�w�6����M�K5�u*Xo�}{O��pQ�!:M���/�!���4����6["�yFA���� <`��m�3����Prr�?���ѱ\t�0�{T��n��$� �(�F!�\rEۿ6��D�n����
]|���~9 ��@^c�6U˅�_����a�u�k�|)1��e#'OD8��~xIYs��N)��ܲ��a���� k�6���g>��m��K=,hB�y�c�-���/����|`-e��T)+�㡑�Յ�A�g\1��u^gX�[18�spZ$����ѣM��k E�9מ���Ѥ�
��f�D[5$�JCDw�mct17�R��^,:�ΊS;�������(%���%MC���0�����vMq\- y�3�N%�Y�40���7{>1(�^�RIo�ۇ�gE�J�p�����$R���:%��;���J8L�b�wgd���wen.K{`(�~@���M�K�8�M3�A�?�'����Tw4�)\ɓ�&� 2��Z��4uqz���� ��"c�A��L���/ M>��p�P�|A�w��j��U.&v� Q�`8���V��V�3�Z��|��ً�vN�{#�?���l��n�S�yz
�}�K�;���t�Y`,^2=;����w~�׶ڛ}�����OZ4�s.���s�!n�(�d�h[��dv�hݗ���Ӵ<�P3���Κ�������a�������3ƾ�8o��$v��;���/aS4�3_\ml����qD��� x]�-!�*�����	�a�ĭ9��7�2�J�+7[���4�k����,��ˎ�9���{�t�=�+~�U�b��Dq���<��H.�ñ/bں�:���S����%Yq�۽4䅔�a�#�� ��	Nk~��8.��*h�	R)DʻGg�j�S ����P�H�h8A���R��[���s��V�e��/L�q�wy�������R���*����Ϩ�/��S�ć��1D�7�e��/1����{B�
M�T�_��c��]p�[
���N�ô� �1%�=S�9�D��T]�.5g�R�ad�a�R�^G�X���;�d���e>��E�#��^oHC���D~���:�#+@����S 9�5��_ d19�a���kjq�ť���c��-A8a���b"Nn�|�|��[y��:��j��Q^�?S��̬j����*B���z�6�D�L.c���m�W�*�:��D�����O�p@S�A�lj��8k��To�:�Y|�!ئQ���������0L[/qP���\�~�y$5Z
�$
YD%ו��r`1��y����`.�-��〪�����HQ�SA�K�נ��D[���L��Ber��h�#�.�ql�Ą�B����~����>�`M���E!��o1�e=���С"׊g���.�h#�K������o/`8q%�\�j3Ei�e�/B��/�G�2��m����=��Y]r/�~�}HY��1ɡ�ꚷ�	r�f-�3��{X���۪]�Eɳ2Ս6*�o���L<ǹL���'�[3Z�0���bޅf�.�g�S�kSx�ٚ��+�s�2������y�S�*�0<㔇����[CSrџ�mHΘ,"��_ǭ�s��T�I�`�9 z���y����4������ؤ���^8@��Ug����3��x�ӕҳ�Лw����"�U�j5�1�%�u�ʰjt�̸;66�
���=~�6�_�(lZ��A/�}H9����M���M���ǌ9>(m�\��ۅ�熨��p�td�`�d��/���|#ib���!jEzx"�^�I�BI2ˢ�\lhk���$a���b[�=�l[�rH���a��s�2����g�Mɤy�QF��y��h�@pMpU�t�Q����v�\�������b%�j߿��B_ݲR�;
jG���K�w�]*��v�@cD{-���#N?���馩�<��<U�Mī�����9��dV)R]�X���������ZL�o4���vs;odr��c<�?SI�"�^����Xc�d��E<�u	xU�_��L��sQ�������dC��DB9���O+����<@ɭ̽8_1��WU�/��9lE�A~�2���=7B_9�e���02��oƾ����KF3s^KGr0~�gK�G*���	�� d ����B�sP��Ի��2�x*�����,s���6?6{3k�E�i�Qu���c�sf�S���eo���3 �m�\>����]����A�!)ˀ���XS���u�Lw.W��	��E��;�U�S�S��H��� 2�jK]��:�H�l{�_J���A`tN�8���./�K#��T�H�F�sE�:�������0�j�/��BNi��������+qO��?�c���`��B�����5�W���Cd�ld=�F_���4"��c���,�(w8�.4��rp��>b�˻�=VCTy������T�גv�l�x����*L/g4x	op�sӎ�/�>�o��g��q4��I��n�������u.���QD�[�* 5�EeӢ�F�H�VXe����*_�܉Ƀ�B�-Joߵj��e�+[�-áH *@O8�W�W3�X�N>Uyu� ��Tx婹_4H�'1:�o�J(�M��G:7c�>bq��v`�B?�Zݔ�Pf�0.�=�r��~2B���]�	B6��:$�8�����F�y���I�_�e�>��pM�+��r�*�Dߠ�%k�_D�m��[]�<��F���Ird�8�9{�3d�]Jkv5L�È��1"1]#~��Ȅ����U�K��R���PjW�9��$6��]���H�>9ȭ�s�
�1+%_(i��-K�����H�r�ju1�G�`!�5u�:.����KbSR�����c�yQ!r%�ڋMrN�͵�WEj�~���mć�g������!bs}��3��P���>��p>@za�LL&᭟�$�e��~�4��v�(x�}��G@���\M�'h���b�z�X7O`n> �@dg�`���<UF�C����޽�$}�0RE��~��+t��(@&\�^�s+U��̨��V/y�Q�w���xEk����=L*H[����9e��n����C�r����09�~�@Ӝ�n���Z,i��)zH�-�"Y_�k��"6uO�ǮNFP9�L��5�[7��uhnp}d1�Nf�>�Rp�{���"s$�=�dt�̟?�Y��2s~>�	�%[�;�������Z�/��uZh�^8�����k�{��m[+�[a/��mv�
1�f�F�!킚T>fp}e�kޏ�>��m�uJ~�D����V����+q�B�Qa��u�Xhz�˒�nu��>J�y��Ư����5V[�Gy�T�\��Gt������+��{�5a��� ��s�I"�<��}�3[�
��sB
e���J��N]O�����~ E!��=D�����g�x����)�t-�ÞMװ46���57�Jē��8��m �R����b�@~P�Ls�\-w�(x�%݆��ʨ�p� b��\ڳ��܄d,V7Y	��M�;r5Y�����)9�d}�0wJC@�$�ƀW�1ef�R��;���ԁ���Q�Ҝf����)}�ښ7D��������]
�p�n���D�*�^1�3���C|j��@�0�[�����n��P���k�-�
�w-i%��	v����170�~oS*W��Y_�n/�T�* 4�mU��Ӱ�-u�sRJ�nLtw͢7���g�b�?�7?,�V������W���;$5]w%
�L:
$� "#��/���1��p��G_�}��Ⱦ���� �թ�3w�6Ԡ� |�̀����x���t���o���돰'�����-��)۞L�c$��>�,)�e�\|8��y�� ����D6���\��@[{�?���;$��U`F4�h�sS�T�l&����0�$L_S�rT]���,��s3��0�Rq�������3&�R]�gÖ���29V���n��%~�k�������i���l� �h��������KE�(02r��u�e��`X&G�}�϶��VOѡ=0��c�l�<.��yT��,lx��Dנ���N�G(�c&��s���v�� 9��N �|�+�72Z�f�`�X�R���bA,c�qB>.\v�3!zj:�"��
v����)Y�e�
�X�<�Ӊ�i> �`M��^0h�iZ��ه�Rڻ��[_�	E>��V�}ڦc�� �����F�y�)߼�
���/X�x:�VBW�3!$�f��m��/�n"�y�e}E�pz�ܜP�ut�_n"(ݨ��c��|!�n�󧨟:uX�0.;��o�'ڨ��#�-��8y\{��[Vѫ��������4�X+s"}Ռ��FMc,�?tO�P�r����2����J�^�!(��m���7��v�gY)���߅O���h(���sUt��������x½�e�$�z~�j=�����J��]	�JL8cjv�ע���O����˪X\�?��:4ʿ���#�#�(�~l��J����<4�a.��$N��u3�9׏�"��=��`�˜Ʊ���T{&��z�&jGm�j�Z	R*H[�n�xj�T}P�ƒ��] d�˿05�`����?ˤ�Z> wHv�W�=�s��s��2%N�&A5X��gސ��D��4eX�^�+]���{���Fv� ��c��1������C�T�
`�¤����W���ޞP:��k�0w(vN?�M�Vwm�G�꽮r6��6���"HS6�ڿZ�8��e]Fᔛ�v�������
j`��̌�?�TeED[�h�n�	hcfaH�����!��p {H��)�Ed�,O��׈�S�pG��l�ؓu��i_y�o4ϕkƶ�[�ډX�N�M�,����?}�vY��8$�(ԇ@�%���[�-���C*q�U��L��T$D����|��՜Q	'������LX�J$dk�=�~��/�{?��v��K�P�
�_���'\�l�@�+X ��g�&�O��֞��	$~>���m;��,��w�Lz�N)ɭ�@��s\�5ȋ�w/�b������&�-G��O[Uh���h�.�n\yDV�p��\^z�ȇ���$ĸ;�9! ªǒ-ˬwv0�b"Pd�Ș�i����ׄ�#�Hǎ�2�aޠ���F��^ ����үBG�d���!���ż��g�Zpr[��t�Rz73��2�����?$mk����5�۽�������mRp41}���_&+a"���R���<��x����h��G��%��h������M��h��5�&�����4����O�67x"��i%% gZb��8i;l����	�����N�\�B����t=��<ǝ(52�3$x�������� *������sw�䑈UJƇ4�"�1��@c���T��x�9����pˎ�K���'�I����0�,|`#�M3�&���&��B�U�v"O�`��dd�h߽�\"E 0��x[�g ���,��Uk�\�����R�вa�J��TI��JC�'Z�����[9��0�B�{hX�j��rJZ) �� ��q�[853�J%�Z����Qx�8�Ҵ��7kֻy����݁�"�զ���!N�n����0�؁7��4s��H�Y"ʯ�$H�
ϒ�Ug�Gd�?���g S��`�8����C�����p�~���f|���<�:��ķRI�#-[�O։��]뇸z�秵e�qz�D�1�N����������0����(2�=��v�ñ�2���-�-�d���	��t�5t��ɟ'���RZ,�| ,?��yZ+�:M'a0��:��	t�CkzG���R�8��MuH�:W�\�s�L��Y�S�����^�'�,�\��hIr�|�
��jA	)= ShWP ̇��~�ײx]~���T�����~�d�cҳ��[��]5 ��h ���TK��U�B( $���M�:�.�~��V����
i�F��X��U�������-RS4��[ߧ�P$�	�Kr[�(q�R�Q��Xڠa*�6��>��z���O�� ���YYl�N.�B�?��7�j�P��kp|�5ǌ�2rǣ���!���+��(-�Ӆ���#�Ț'����ԬW`jD��u<6�@�g� �皝�%��k��_�۱�9����
+%��6:�jho^t�61k'4>1A�]I�/�R�|�+ӎy��YQ_���QQWaf��T!����U4�if�[C�c�2�O��C":N+�w���uP��z(�X��<��V�����6+iRy|3�2�D��L�[a"_���u��w�|��ʩ(U��2�yq)�(��}b	 ����2��Ϣ�?Cԅ��3ؿ�ؙ�;�^&*�$���9����&��JP��Q|��ȢO����Woqy&�>g�1K����Kf��L9�8&/0��Qٌ<�,��%�3�Cg%�6I#����G��"��(O/���5C�R�d��+.q��eih�W�sx\��|���c
�c �R�L%YHy_��C��>{����bF��5�~�u��b&��{�8:P(ySt�y���%�P1AJ�n)�oP�=��N�@08��q`k���"z,n��LSU:�?Z��w[�81���L�4��ZC��h͸�:����q~ॸ�p���l0���p�`̋u|�V�����t,����nR�;��ձo�Ĉ�A�Ef�ҾND��Ӳ�@:��ނ>�U���B��0{���L�`�/9���O^m�H��SUY������tR �yїj]:}1f�M+y�pU�0�H�%o���P�}ũ�yp3K�~�0���q`"C݈����i�7��|:��F`���;��v]�ƌ�TQ�������"�m��g��щ_�3$�vbw����r�cXe۟����ƙ��3= ��0̤2�d�=dqHXs��֋�~sB�~5e/��^�����"Rz]`���ˍ���])t6R�{��?V��yE���Z�֔F��F��A�\w��o7X	@��5�V�o=Az�	�����wi���$$��H��͑�ȱ�t����*����mY<������wI�	wY�wiEJ�c=�"��,q���U l_ŃI��Aף/_�/kG�9�`���^��4)����f�%+�7��Ye6M~�J�*ǎj%���'r�p����GR3k2�Ču���o�O�;KE��O�H�爐��0��qs�N��×I��͙�^(�ͅ�[�$�Eb��7����2P+S��(ϧm�y;�?¬9��E�dU��<�����,A��_������G��1�~���(~@�]�^w�'�P nZ�W����s�l�K�RNֶM>:׀˥ �� �Q��R�2��զξm���(�*"PɏhnU>��6��)rĩ����>�%	�g��\���И�WQ�ܚ�h�-L'{�%dG�@&�}��gy�w��i2�Q��X8*-`�]��\�7����M�@y���l2,���j��^W��s���T$YPty�[F��8�$� g�����F��?t���Z�*u�AW��%���R;q-��P�o���tp;8V�(���o���]5$�p#Ё�4��0ʈ�qJ&DE�NMCd�hC��xe�"�����O�Se����i#־s�ǥhANq�������d���[%/�rs�d2`g��|u�K�ro����b�2�^2�A���|�:wT����1ǂ���z�`��n�Ԙb�Ǹo��	�3x�@]5�Q�>Py(�N�u%I\�>b-fQ�&�y�<3C�F�Zi���,�l�,�)�h�;fA���E7y��z<�j��d��u9pd�?S� V���	S�R�ua�EƜK_�@����g_�.{�x m��9vC��D�M�ܶ��z%}��Z�@}#�z�(o�t*,i��1*�N�*�0'��Ա}^�)����[��ao�d~��,���z>��A
1����OPD;!�פc�a(�c��4����.KS64=���2MO̕�_�*�-D��:H��f��(�z1'��6����\x��40��`wI`�o��-Z#v�F��[�L��U��WJ����-x��>��
V5������1,�\ l�9�6��� 䣲!�\�+��2��B�������XQ�)W��F���sÍ�*�P���ʂE��y�a�dͤ���dOT㬥����Ƶ��5����Hr	�u��"����50��QUY�l���e��ZW֯�g�U�.=l������6�
��k1������'	lFߒ#GjP=�Tf��%i�`:a����.no�i[	|'���5��`���P�J��h�{���6���"a�\V��2xS&d?
�LtU#8�ln�-��|�߻ ���u����B�:J=j��M����rA�IU��
P>p|���ȃ�ޛ�h\^�99PX�a1�_S�����5a=*mx���P%�ӌ�n[�B�+&�2��F�l%	���K�:4d}���H���7���2����C�LBs. ѡ��-��/������mg�V7Rm���L5��)?� 2S5*ǨdU���ȟ�-q�q���D!<������0�Jh�;Ble�cj3i��u�b�s*C�K�``�}��@^79+���"u��Jjp&���AsF���~8\�q(}g(iCP�������u��Z�i�CgQ�\�D(m)f|���p��)`�K��qZ�E>Jr�)"AQu�.�*]�g�B�Y%$	W,|dUs�V<Qk�h3s5z;^��|A�� #��n�<{���@�#�;0�,��o���쑲/m��2��Kn[��m�F�x��3��vT���Ur��#"�a��z�m��'�=������x��6�	�6xSv�,��/� �j�Y�Y����~���U8S}J(H�G<� '-	���'���
�Wk��� 
��@]�6�������1��y������a-����-ڮnrD��"���	��C�缐�~ǈG�������T(SL��[R��<B��5����g����h[U3����]�v�*u�̡w#Jp�7>=��j�X�O�\,�{=�M�����d���e0ݰ��J��:.���Ձ���M_����:�R����D��贾x�Z��4�t}-'l
z��U�rR���r@�/K�:|��?��K��ZV0��L�]%8h[�TQ��YX�vx=��%D8ϗ�J&����=ͧ�ݱ1��:zH	ܞ�V�d�g�6�g��п�3��mѶ���!��,�`o�"n>��i�vf"��H��<_?��r���W%vl5sQ�c��:H���1�G��gW$Lm/mIg�֚��ʇ�]c8	���@T�L�s��a��Ձ��Zo���b�?����<��iz�|O��6vWbX��䩛 i_��9�x�=�����Ŀx_W��ߺs��i�V�X�9�X9�zB�02[39QO�[HGSbyi�Y�,$'�� �w��m��U�_@c�CƷ�&�/��'�����)X�@4k�[�4&H�13Ϸ��|y�Q;siF簺4��]�kbj�[��yD/�x�>� f�3��6�6�V������nr�7�ǒyJ��%�䆉^�/��{�_�
Oj�L�.0�$w�*z�iR��O�9|�x���O"��$�2>�2	�#�/=m >��n�	,~� i������� �)�h5'�Maի�_�-�a4���U��$6���nr�ߤ��lP�Gdʨ����UZ�N�.������Wx�$`�������3n?
�	��9w҂
o�;\kO j��g
���j:̜{3G���C:@�IDF��9�"ql�c�ި '�uHB4�=�T��"rc8���uE���C���V@0��R�r��v�����#>L�S���zA�WJyă+%���[�����b�z�/�օ����7������3Sy�l�|�$���N�����qw0�B��:�/��\�����uݱ�_ٍ���D�s�K�]!�	�7�"J+1L�i4��O��W����AR֙���^g�+����'���Q�Q�����h���+x��[O��DhPX���h�Q�(I�"n��2�F����l��ÒvuИ`��:G�^g83�Q��s�K����gN�u"�ɗ����K���DeL�P�p����g��,�+�����9A�iC{�O���<@h�����	vX
h��0�v�\$��5Cd%T[��$.[��aѪ��m�5��L�ES�J���
bk�ƫ�
^���̵_�n`�i=�������Bc��[.@�l���E۾�9H5ߙ��7q$�)F�"慗0�)� N �+ �mS>��ƕr>�~��w�X�SϙO��X��.�Ö]��Ω�ғ��_Bf��f�n��0��R��u�"�b���j;wYb6N�K�e�J��SR<h���ߦ��b�r���Oh�H��Gfh��
�zD̊ �i�a/�́}NՐ�Nyy�i�M��U��K� !��@R��}Y��9����׈�H��n�Y�췾�9�ŤD���o*x�N�m3۹����m-v�e������K�=tHZz�W�U@�C�B7vo\���B}QWb�l�ӥ��@~��׈@�xK+ e^����A%�!`ƍ����z0t��W�/�Ʈ���*�t8�֐(��bkk��ԫ���'���]'�,�]�W����A�s�)�P45�p�!�a�Y�09���m%��g�H���C�'��\�P���2�G�����27�D�rR�O��"Zh�?Y�1��"l����uL�5Lf_J��|zyτ~lH�����k�5��I~�~����%<2(��[<b�&�ழ&�Mo�	;؊*hΨ����kw"��ޭM"����q�q�;(��ֿ��[����6:��p��3��'-�r�@@��,�R��O*�[g�Q�E�oE�����w�q��������R�e����&�;�D
��Tk2�~i ��"Xs�0k>!��[40���b�l<A��a�Be�a[[�{��5���5ٳz��;Bx�}�w��v2�퍳L���~�Ɓ�tq?�&V,����d������Ã��m!�;����O������G"w���Z��T�+ܰyp�i¶���g�;��~��m�1��Y9�T��f�0�c/kO����+�ނ	<��@d��wI�)	��Cn���K�JC�=-����q|?�f�_)z�侯����LIٝ�=a�<9q�d����������s�اj�-�W�7�	��S��2M��aVR��p�q�~���N_���w���R������5�#?�Q]>i E
��ŵ�ތ7������u�����}����u��2:'0�R�-�����.�8�%�R����6}"�Q�9�C�͏�H8�mV���0Q�d�̧ų���歨�닃��1m�$0��{��h�����lr��:���!KD��.���\Kq#��&�S0i\wt#U;��4�����k�S��a��V��cǝ�D�1(�Qp�t����a_
.��,��̵�3V��q�P⇈�)a�n f1h��koZ�84�x^������1 ��l1��c����?�C��]������$U�jJ4|��J�Y�'������@��c�M*�cZ9봩��/�?�U?{�K1�;A�a0X�nA�(3w��<sxrlL��n��!WS}�ZC�<G�dv����Ν��J-5 p؇�:[H�Cm�DlZ�����YZ���^��e��>�����(�ي�e��8��r�9� ^����A�6G�tu�Ѧ��l4I�����z� O�v�}֣�GU`�i�G�`vX?~S4	�v��=�T�{�n>_D�V���f����R2a�|6�5@��:�!���U�Z�9����48��ƞU�A.������F�Y����Y��7|��-n��I�C1������	�������Wг�\XY5��0AUE��� �_'v�FG��������-��s9%���]�mWq�%܍ڠ~����&��o"ǜ��j�с�D�
<Œx�]�tU�~ס�%�v�Ms���.�U�:I�	@��}$ǎL)���5K�����"��iQ�ǣ1og��jeo��� ��q��5���8&U��M��O�Rۼ���+���,�Y���N���� u"fS���h�T�\y����W��p����Y���~���+^��%����������b`y\FHc���%0���+BG�����1J#�Lw����y�Ҍ�.�CB5G-i��w6��c8qIE�־p_�L��P�Tl\��K�>풯���asx3�V�W�tH�����d�n���Q�G�AE�ˇ�rս��zn��ɏ�5��X[�T�ci�W��Ѧ]�*�����tV	��dFWd*
��YI%�Ò'���p�gҔ�ڔq<
�I�[��%��a�|�Pk�>F�:.���t�6��c�[y���!�J�\�'���襢t��Jr���l���r�k3�Q�;��?��GQ�ŀ�"v�i4q1e��J"3�y5�G�σaq� Pt"�R.�Uη��(�"�z�ˤ�T���I�,�F���lg�hǚ(	�?��{�|/��R$5��ʹx�T�9{���C��i��{BO-ʧa��Y!RO�m�j��P�CvXRT��A�=��.s�I9�r�a�u2�O<�/�K&�K�������d�hNDv����2c����P%�4�W�ᙖ����(dH��f�3�_��&���A�?���Gu��v{�9C���7!V�h.�ě�����ce[}��!�9.����P/'�)����A�1"`��T����-�߉ˇ!�ZF&�'�Ay�58l�Dߍ�Zs8�F���rq[2� ���C���>��'�r9�%��ՖDG��	�*�_�Uu6���%?��F��~����a�	#�AQ��g�� �S�M���~��F'�)cx�V*��#��<�a��y�,�〇vnU?�z�d�*h��曃 ������L_	Yd��;��QP�#g3���ô�둺Ǭt����&[�؛�����I�r툧�y$���ĸ��p����^	�U�hV��}c��WU�yb�/Gr��ؖ�B�r�͞�9��N���Y߯Xn��*
Y��6�MHP�2�_dUV\�"yG���%��զ栯7�
#�bM��Q-��D���ǫj�R�h��Os�4�Yqkd�X\y�q��q��C"*
{ds9BI�ql8�A�Y{Yhcuo����
�1�C�]�r�$����\v�nBлK��v�\�����~�i�����-�Y�&^,�"������Ɇ#��JY��V��E�0 Mf@3��/�ю���]Q&��X�}6�~_wB�I��	�)|���� ?*�l����� C���x0M@y���U�1��3QkߟI�r�O��RH��5�,���ʅ�8ka�~�u5Xn"�]N��Hp���pj��PpbB0����d�W�p��9�Ҫ���$LlSD�U٭�ʥ������:���Ƀ cz/h��aV�-�c�A��[������in���b�cz>�A����Υ���%Jv;���a<�@�����ƃ��@s��M$���]�Pz�кOB'��)Πr��`C��n�Wl��F�wH�(XtW���9u�6y�y�x7��T�i�8�w���͊u��9;2;K��Q׸Q��H��	8Yz�j�n�jF�@�ƣ:�YG^�\5\-�+����:�٣O�:Q�/�G`5D^p���5�m�k��]�L8�E d0;������G���t�޾@��EZ���~����c:c�(�lL\ ����5��3wP����W��Q�
�=C��"��������l#a����^<ũ�=����ב�g�����?�pF[����-ak
DDO�%x�30� ��סt�������OB�TP�L�h'il���g��Aq��#�&I��{k!C_%T�'q�E.��t1��_��#��}��#M�J���ߚ���e��|u��ϭ�P��,NC�rߊd���r)R��x������3,�~���+ц6�3���\�U����''h��,�����sK��U՗�}t|����XB�V�^��p��S�a.��H)��ԼtQ�Y�������Z_�����ϊ���SƤ��A��z{�6�Z���ļ��6�{~�!7LL$�����3�#��q���������t0��c|�B�6�����7�t4H��=�q�C��&y����_e�B�ce&���<
�1R�O%s��)���T���$eJ�QT-Lv������!�}�I>�X؂���L�=�BOuxo�dԿ���D��|������7���y:U�y�IOׁƈ�@���r���v��NAb$��U�"���O�!s��C����JSf���r&O��[RZǃ�����i�8� 8���0��bP��؂��7ݴ2IZ�-����lI�G���^�1��_t����d�(�[�
��qfg�� bm����������6MP�A���(i,de��Qu���]c:N�4�;GY>
��� &Ҹ�e��NB����'��멙N.]�Wg}�Z�H���3z\�B���4����s���RU�V�����9h�_7'Ѭ���أS�����B��4������}��{�ßvi�(;�A�S�mtPX���>��f�3pԌ���"Z)
�����@�9���tBт7�C^��L���_����T��:�]5�E}_��s7��	2&�7Q��]|1�Nظo���+�~�����ɗV��3��Q��D��.`q���
=yXg̱�jC^M|�]��HF�+�DM�dx颍�z��|�eiemoJ�|͒ij�9��zc��j�W�{&���rHpA��C@��:�h�J��w�v�(oX�|1d��[&JQ,ǝ�X���4��D��/��:{�}�D�xt��U3�V�m+���i�Ժz�MX�M��Eۢ�A)[�?����Fjt��b��J�;R�MM�^��!�=Ũ%E:ݍ�>c5����F�{F&g��6m��_mh! ��p�~3I�Y�=ղ1�/��R�'�"��|C[Y:ؘ��	n��b=�����{���`G��>Կ�ǂ��p�&\�vd�՞)�?U'��)vp��a
��2sM�������R�t�:.��2I\hv�6AРgZw\]�=v�f�����A���n�2g�Ds��:,�_xY~�v�v���E�f[m%�	"�(�y���(�2�U�'�����C+���)�L���F�%�Ε<�E�L�P1�y`֪���0���J�;g	����k����GAc{��l�vc��JM��Q�c�hfAU�U�D��9��m����|K���q�9��Q�$PMS����jS��b��J�P�����Î�+!,^n{@�GY\m`-�qw����g#pb��}�|A�6�»{V�
lɨ��BE%�TR~Q�i���=T!Z[�F�'Q3�%�W�R�ŌL����Sb�Ѷ�&1�]�&�w�(�Q�,�%��O�N�!nĻ�;�cM�V�?Y��ʔ�4�c��V�(��B<+&�I�ܦ��LTz�f֘sg�`}S�[�)U��1�	:�'?��+K>!ݑ�m��oos��ܴ�8�J)|�6��<̏66��D՝Z �+�)�f���j��䋂m@%9��6T�S
mNt�z��'i��4��K��(�hQ���s�^@?�	m�ly
��/�~����G;5o��Q���iN>��D�Wc�WR���2M��-ه���&hI�k�����G�Q�Z��Ld��|�I�djGz�k+Ϸ�%����E�a��W�uӋ�E �хDY�4�e������� ��L��H��.��8p����3~vA:�y��aQ�J_~��/: �t#l�dR.I�4�/��r���g!�û�U)<ѹ�IJC
t�p��3��_�"�ό��PIR^���7��������Q	��F<�un^ɧﰈ�����c�҅�ZUA��;�?j�0���0���D�x�]��XX�.�&�5w-�UT<[v]�O���&����*�!ݒ�[TP����9��o� Y	2���c~��>'��J
Ŭvv�Z>nِ\$lrL��y���Š�Q���4(/V�0]Μҹ�ֶ�#7g�_6ĉ�g�{+e��+���f��*��(�_��Y~�1�'�(w ������'q-'sv��ը��f� G����jі�w���F|�
�b�<�D�z��$]2��b�y�j~��� B~���Čڿ����B[�˪�N��9q�����U�z0C�.J�F��qg�B�;�ԉ`� �T���\����d�@�S7>�0Y|߳݁Ɖ$W��#��As��.�tm�"�U�Š��։�N����Z�N�����S��ijJF�vQVWi?R��H?4xI�℅!Ec�; ��s�T'�i����ь_*�n���r5�qc̦`D�\3gl��D�?�+�-�}�gr*��ۚ�¸^�u�6k�!$l���P=�!L�7�\���/����{��T����d��+:�+���;�î� �0#Pt�����EJ%�Ir���ل�fV��\p\ګ>x���Sɺe�1%�(G��lSMSz9�-����g�4�����W�`}2�ɯ���E(X
?=�5<���_�Ńd�!�i�	:l�����P}�=d/[y�}j���9�Ly	$2���ِf������e����?�(�76�!c��$^��)�U`��a&���hO9Kv��c�P��mI��=".w�D�i>{��)�t\ۙJ���ѫbS�	� �T���jm~�ku��yEt�,}�$�oE�Tz�(��^L�K��ŖC�l���*���6��4h�I�ٺ��)O�V8~�*�c`p�(�dVШ�nJ����h��>5P�k�����7�_B�X�jd�Բ|��W�	g~�H�)�gʬ^��W����|+��Ǽ �DF��u���~�
q������أ%M�'�9���G���	N%���#J!$g�V�j���2��mg��T�8�<�Fy*ּ����C$\(��x�3�2�(�����5��-�v�O��g'�t�Ĝ$�S���B�K��V��ҵ��Dt:yeA�Te�SF='��	�'��ʅ(��e�m�s��ϔ�/%�k  OLQ#���o�'�N����w1��[)V�p�]n���S-��-�!�Dy�1��!N�۷n�� �C�Y�z3�w�'���?JSq�Bh-"���V@���)µQ�:��j���<�(�� Ʈ�4U���U�s�gSm���x�YB���҅�J����;6�g�61�\~��=�L�6#al���Ѧ��nV�e�R|A�
N�.�ȿ:�X/���^6�ft`b%J�B����9�KU�g�`yf�?���b*w�uǂ�\�D�bŻ"��&Pgҫ���"�G��D��!l��w�A΀�21�S/�(%��`��u+~Zr���4?}� {y��/ͻߴ/P62t��Py<85-"#��4��s�45d�2�P������!Fz���ۓ{2_�.I�3�z{�$n���^C����8|��f�7����ؒq:|9�P=k�TGh�΁�ޛv��]��0Gs�;'#4���~"ޡ�I좋�6�d�kZ�c6?Ju��ݾ�����l2:0$ZLd�4li����u!T s�$�|yqR�:7��'Q�,�D��6/��L|�vrJ��p�q�TBx�i�ǳa`f<��d��BE ;)8�Qʡ��^=��_���T�8cc��D|��Z�ʈ�,�cq����۷a��f�߾с��<�t߽n7�˻`M˰��fWN�}Ek]Urk��כ�G�V�$.���>r.���e���^W�o2`p��U�\�zp�aӰ+�{�L��0X�U�J���I2D�\V�J�N��y�In|0�@Ǒ ]�\�з9Ay�f�ϻc�'0U��X+����ZU���|�� ��jg�!e�������6���	M�;1s�Q�1�v�X�+(�x�!\��A�<@�s�Ba��g?Tc����&�w�c%���ken�NhՋ{!?�� n�#T�6�Q��iz�5-� B����
E`�1��-(�B��N���5�+�zO)���P�!�A c~҂D~ [qjͫ;S�E�]_n���ϱ	S8V�zB���S�,c� �t�@��6���Ah������#����5�(NU�<���j�>p��G�~3�����^�*�1U� ��l="�wQ�L��W��5���5���yz������P�܂Q��v����IߑT,Bh��5I"Ϭ�3�_����8a}VBCū��s+E_ʦz��2�9������M�wj-��G����S�z�W�@��b,�L0b�|GAi�� �#&��B�nҭ�:u��/$(s=&|k�����8��������2�`��Ro����`��*������l��΁�LV\�U;uo;8[���Lп��d��k������LlCJ��Ny���|���e�cIu�>�ĳ$_�ER5O����ep�n܀�����fl��-� ���}�R*nI��^�-�;���~}�F�~d�M2�Օ���\b��J���cJ������D�}`���Ԛ�n��OvZ��_ (�S1jGo��oMgm��<w�_T^�T_�{x2�b"͹u0[Q��@?�i��6;㯊�(i$m��}�����V�<�;M���|��\�R���@�J�{��nXV7J]����^Dѣ�V���fe?�3���J���{[�{J�2%>���%�F��e}���������O��"�>�i���**��eB�� �B�/#>^�v���+x�ņ6%�o���Z�+����+x
��4�v���8��s9T�o���Re�I˻?\����$� �E+���q'�p`N7nZ�ѵ��.�lU�7�g��C�Nn(�)�9!{��g�Ʌr�� m��\l�7��(~�qz'����O�$>?Lso���ڸS�]4���1ŎSSD]��	��HĈ�07_�Ǉ�oe�&. �v�b��CL��Y��$��Եm���%K�}i�2�)/լ:ܬa�=/7:��hP�O��E��8]�"�p�k��Q��d����̲�����.(� ��O>�]�tv�]muK��Keg.U�n)s���ޢ��1̭��WP���2�V ���;����@�,�� �j��!�"`K��4�g@(Q�,W�D���(hm�����"&ǌ%
�F���"����������8y���vAEk���աR}KA��1��a���/�(ج1��S��o���l�cvr>S�� [��;��x픩�����Ƭ�!����?Ⱀ�)����ɑ�=��n���K���J�#@�>I�C���1D������]5��Y��56z��k�����$�x�Z�O�M���N4W@?��"�k��#��%7FK_r������;���Z���a'�JǊ��U�J�������e^ԥ��2丣a�]��\*��d��R>3�Kg�Z�3�h��@�^&G}!��g��G�}E1J����~��"!TJ%)��XCM�lߎp'��R0Ҳ�?�d�0��=j�~v����i�~[p�t�~��r 5����z�h�(���4�H�y��f�P�l��� D�o�C?��	�d�@�vct �TxRk��ύ�I9�
�n�{+�ޤ����q'�PN�KTk�n�0�6D�_���<�p:)�rwy6uJ��w��͆ܶ��P�]JG�U�PM���$Sy'ǥ�IAe���om�B�3O�.[�؋��%h���5'��O�9�p�y�cF�7õK�6��H��D�m�!�WQ�E=�����/l$�!�;�ލ�rW��/M�a��/���!*�4���$�Qrx0� �pM*��2C�Ί�ȸR�j�=��
���	異�-?[D�	��g�{���}��78.ⳃ.)���o�����s��j�K	��X��ٟPV��~�L�j�r�J@��T1���sR�I�^����H��f<]��Kn��(~gmKW�jZ���p����t�Q��:�$	�{w��'�*�㮳Z��<T�-���y�9Ҥ�s
�"� 20��P-$��u 3 �	��A6� G�TG��j	3$��*F#
����w�ӳl̶�h8Z��=�c+�t��ӣͿ��\��A׎��\c�#US�šR�顆2 ��Ұ�^E:W�%���ĮP����!`d��!}�!��~���S�|/ug덋�y�i4�Ļ��Q���Ai�(/_%!�i'�df-�����A4�k-����"�А?Q{'K5ͫ�K���W;dS��]r�.əB�'yr���al�=�>]�Z��U�1;�A������8����
���|���hs{9]��T�ی�
�WN� I�k�uٺ%b׏7��	�� �m��z�כq)^�F�Z�?W�IoR�Ķ��t{�O�>�^�L��xt<�HdS�T�	�%��N2T�1�o|�F/�Ȏ� �	W$�w`6k�s����0G$�Y�f��]�O�Y^d���`SS����=tV Mߟ���֫�׉���{�rM�ZQ���E ~鑁�rW��
p������n�:P|��GI=ӿ(7��V�!ĝ��9���0}E��8%)�(F�n�XY{�KbӖY�[-'֟�}	n��7��2BJFcb�.�v;�yRѣ�R� ��o}���OW�e�#�G�-9�1�f��'Ce�q�,"�od��r�ۦ ��?�hቦ� �o�m�l��:�e#('��~�L���?�ELCO�Ȼ����}�C��y�9QM�8���(_
��̩���N�t\:v�^�}�?9�^B� l��߃c����ƙ�l U��]���3�&�)|nGc���1}�U3hZ�i-�g����8�f��;��C"w� �r��"�0i-;�(�T��Hkpтݎh��.��S��7Z���JCA�m�hz�5�T�PFr	Ҿb=︡�H+�h�E��O�8�كr�f�&ʒ%]ߐ���+ٺ]�?��O�\ٸ7s�R�����Ux��k��ã��־(���#(��`�#F�76��[-|��-���5�
w633>S0A�x81[Yp]��L�}�G�*��z�d�#ƧR��LZ��.�q[U���V�� *���>�oB�:sߑ׬��{�߅�m�Mgy�,�צxՍ���0��3٨C]�+}˞�$���#G��;*M�:T{�Ȣ^����ǽ�L9l��-P��ژwX�&`L�Y)^ΕiE-�l��ϟ
"ʷ�9��me���J��Q�Dr|���5<A�D#��Խ@T��#j�~pOuxv��	`�
������� �k��?9,X�'Uv0�C��ZD?$[��q\���
���blP�t��|��7�`,g4t^*�
U�BIW�c!�5��]��O���;+EBP}w#At�R��&Xp��*�� D l�OCgn�=簀�sϛx�z����w�)���Lbo3{K2-Ҁ�f&���I�h��Te�Mv�/���M���=�{�F�M2%zM�'"w����t^6�� a���+\�'1�"i���6�o�Δz�����1�S�P��h���@cR�kw��>�J�Ē��1����f�#WS��-:.T��#��>���M�:�N3�h#:�!��A؛�r�;�������}!
���u ��+��[���pؼ8�|!��=��W	|윰�装d�qT�H� C*�� h�UE(�@CHR�����Ś���\(o�_|5I���Z�a�H�G���9��� X��Q��c�SGlL7�5���mOѬ!�?iՅs)�^��o��h����sia�����Č4t�F���4�-�)τ���x������o��4��y����'}:r _��0���H��0 rsѰ8yuQޠ��`��������sn�+��J$�������Lh���P��p�I�X��Z&��ߣ� 6*�<��O��~�Ba��@�&���r����;༶ިK(��j{�Dc�=~/�Q�q�Ued��o�Й����̀�HKۖߤ�	f�4��T�#!���
����1nW��辰a�[�%2�.����C��V�,n�Sp	��7_zT�� �]<䤾����\J�W�.@c��[j͆�
���	�O5�
,��V4���ƙ��VsaĆ�MM���1��&��q�N�AU��I��[`%bWb�5��\��s�|�0�*/z�Ħ�Qc{����m��y������R�̷,�I�5��M���i�1�;o���Di<��;�E��W-=����Fң������<�4�������*�ΊhOh� S@��nj��b�~��R��t)]��Ck�5�G����ynۉ����n�� ����o��{)<�
�	�t2�y�Y""g3雮��J	=u�k;a�r��ӕ�C&to��M��Cb��J�2J�(yy!o��Y��@7܄��̾(�Bk��������h@P�+zT��](NY{�)�rky�!�O�N��~�k��l�K.��Nd�������_ЃO�׉�<�_��q��Sų`��i�d4h�N��+i�D5�J�u1XМ���P�ip�m1����[���g�b�2*��-����l%7V�ԲV\G��Ȫ�Ц�ۇs�ƻ���%�:��$4rh�a����7��3�Ŗ�w��ǯ��B�Rű�pB�"f�s��^jL�%�9�l�_�9��p��p���MrC;�ċ������}V���\QZ5����?��R��k*������K$�.3��m�M�n]��<��;��@L��%�BW�\�݄C���*�Ʉ��1%�}*{#o6�tlx6����S=�%*ՙߪ+G��@��)�Z�\�z9�S�9ә#q��C�V�CN.��v�فY`S�(�q��ua�,[U�C�۫�>[{S��1�j��4lھ���L�D��7���.��\@K*�ι��T�	H��'���gC�wn�J.�rd�^�6�(��'� �V���˳M}�?۶�;7l�8�:���sD������Ʃ�K��h�^�DC7Ld���2� Q	�� r[����̓� P�|O����h����@Y,�O��1bv��}��-��pǞ�(J;��F��~xG��'�() �
 �"w�6��C@�E��X�Smz��q06B;Ƿ��^f�x����6���8����lBp0�_^I�,�8Y~r=��*M��ki+�h�v���[r��Wu��J��7�E2V`~����T��^x�)7,���M���W�^Qs��P[JP?6���:��\��Lz�'|2>�~������� M��/�
C�J������/)�\��8�q��pǔ]'#���ՙ%�ˠu�'�  &�bv|�X	�L���7G�d�\.�O�p
�L��Q� �ޙiך�eO��`v����s��i�px���]���Lf�:��'���,�)qs&0�U�L�kV@�itw����?1#Q�K�$�S�T��,�`k�٤vJ���@
q ~��W����T"J��Ƙ��D�G􁸠]�K�Ͳػ-�J�AFZk����C����V�+s�o0W���
��H�n�G���2&�XJ0�����ߦ�k�f)���Fr� �wx�H�X}H��42�,��O�f*ly������N�r��	z�s�r�HK�#��qۜ�g����T�����Kę�>ъr��Ѫ��nȎ����2�u� �
���Ȑ�$�Q���uV�Iv��_,��xV�Б؝>㕒t�[�i��X`R{ג�/��u"��L# 	<ꐰw���--
�}>�o�H�-2v,铣֝�cl~�ES9(�`�n��2�WP{��g�A|����o(�c�ɿ_� ����8&z��0 �
Yzk��5=PK2�`��9�2��߬��أ6
Q���Z��K�N&�H�g'>�I�Cb��J���} 33��� �W�>�rq �aԔy&�k�m/%�i�/C�
Z�5�49�S)OGN[�b&^��p2�C��������7�Z��qO��m�q���Zd��
(��ZO��B
yS����G�c�����?�m�٬�3aM������V����΍	��s+�Z��6al�kL;I5(�Z�Bz� "���lt&�]"^.sW�ƅ�{�h������\�*�d�ݠ,����0���"=lS(��k��n8�����t�]9�)����|ސ��O̵e@��^�0�đ �w�Vn���ޥ��X�M�	��4YǼ��-�f��de�0|B�R2� ���baq\���T���E3d|��Z��}!N��~ T����fQ7@�O7��=\+sW  ��
?}�X	���6>}�%)U�QV=�C�C�����DTU��Ҩ^q��KȂ|���ږ[�5�T�(���ocu�]h����M۲Vg�	G������;P�C��G2�09��o����L,÷=,�J:6��ҫ�*�{O6�/�8N0ZJ���6�1���{\K����1Z@�FDK푰��?�	�[��Q�`h���T���R��c%��xے��d�G����O��)0�%�WzSI��p�G-	 ��=�X<I$�񑋆9�E|-��J=�\�\���k2	�U[�{��_�GC����E�0�����<9��3?��֩���l�t��=�=�$��U��-j���j�D���j�{��O�7�'�j�ᜣ<�v�Y�ܽX1L�Y��vsV��R&~�@����n)a��a���RM�qڱ�T��,?���m@K�<uG�ғ#��3*H��W���1�*���^V~&V�������'O�I���d�鐰�jf��r�c ���ھ����H]QwCN�_g)v�5�!^�s�n��u�p3�����fo¦	>�{!�J�����7�4�kg�*c�Œn�\��L�ڗ��a��l5n��
cU�N�>��l�B���2��P��Vg��ރh��0��%�o�5=?}<���x��N�q0�hȠ�+����r�%N,�%6n��m$��E|�t��k�����[N�
��T��{o�F]��p>X��H@u��HU9��z@;�{��4��P-}���ϝ*�u��ߖ��i��?�|�z}Ȍ�-����~��}s-l��c�4u���贴P`,�<�7"�m��s|в?Ю��6��6}���=kGt��7�oQ���wC�7��^�Y��q��) [U�*p�0B/wTV�~DY��*G�cܙM�Z�
`䋢��=	��]�vc�ښ_��Y3t ���dg�J�����e�8uQ��@���]�Ū�k {�e�XV*�p����&�?p>t�Rc�A�!&k�jU�tLQ�v�ɼT�%=6ۜ�/h�ߠw�5M�[�tX�U�"����õ����W^�A�垺�0�R05���}($�9��d_]Oſ�v2��vLMG|�1�T�� t�}���z�"�+�YC�ǐcXV��_}y̯��|�[j�w܁-��ޏ���D�T�>�p2��^7ࢤ<B������<fľ:�AȚ51c[����)j�w�� �"V��X���F�,τ0`�S�s�Zwn(I��U�����Y��Wt�AGf�<��9��vM��b��`uՓzA�9ŭ��|uGN�?T��}�9���}{���w�%� G��SN�Y� $� '9:F�b��K�nZGŢ��;�T敹V|���8�:u�nnj\�(3�/'�_�KS:ڄ��@�Al��I�pѸ2i�'\��s9c�'w�9g	Φ�x`�F�5�֭;1F�L�]���i��z��-u#��s?� {4��6��0mN��;���啚�i��?��E�hzcKt�[�
[�e=�P3΃q2�	�S���I�z�~E�PL� 2�b��W����}��S�5�S��N���λ���O������!f�*���]K_ϗz\���@t��>�KR�!������O��R��nd����0\~B h���!�5����0�������
h{/�D����|K�s}�`+|�S���P޸!&ݶ"����7�'u��&�[�?m��N��$������=�9�	�1ܬ��ؙI)Ȋ��Wf��hJ�P8�09~�GgV������8ӷd�H��n�����
'�1Swtݺ��dY� �����2���������G��_���<΋漂�pn7���
Qz{�P�V�?n�l��)��Ց��c�7�?7?�����b��|�$`�3ʾ)����H�"B*�1K�r��3p�˩[/4��n"&R��$�,��<BmW]R�(��$M��sM5�yN�j� bY�ͺO��h}��%��J����_�}�)P_~-��H��X�i��USg�&L��X[��僛W7�LU��s��#��O��< ����܈=�?�F}5GI����u��Ec�F��m ���KOC�n[���'>���y�	�v}5�_,1gx�	�w���Й�ɋ@����N��<M�������݉�\Q�0-Ӽl��q �[�@�����c�vJ��C�z�_ح�q�y���J�_%u&a1�B8��	�I^��jZ�%^arە�w"\�����nN��;�\D؏�l��0�pt���'_��6�.F�A��$?ӭe�&��uw�\�6K)D���|�O�������˘!'�yu��EKL7|�?�p��v�F~P��ސ���<"o��E����G~]�B���AQt�3ud��3���� �3��q��d_��}C*e��ͻp��:�+Ό#��Wv��y���\+��(�����M����(gs��0�1����g��@D������|`\��3.ٝ�j�YA}���qX�c�=��/������&"ǣi� z�%҉~M9�L�R�*��l�9׭$�1X�e�p൉[�M��n�z?�n�wk�T�W+��d��� a����Y��MXn���d��cl�oxYAbZcx���&��2��a1�{�>�O*<+��AU���Vy}4e�H�W�vJ��^��:_�ۚqA=��
C��'*�7x���H�����zLs?�J_mz�2'zO��P;%�8�N�Ez��ȿi.��z�+gbr�`��)N��'�b�X_���꥿".ޝ���.x:+K�ǲ�n��$6m��@򜘹����Sc�~����0W' |�q7�}Z��/���t���N4_��4��uƢ���$b��[��4��3yc���]N���Л��]��C�hU��W��C̓S^���>~b���^���yn���<��q�� ��`�E:["���$rn7'4��/|%w��¼Rzd���	�l� �=��+�����8j/��Z/W,۷0��r��qV�v��tՉ�v�a?��W^!���W*�Ǵ�X�` �D��ͦ����$���k�כ��:�.n�j4���w�E�����R�[������Q���ĴV� ^�3L�\���~��{� �T�3�p4��9P�RXl^	i��e��n��@A]cV����\x��4UTYJjQNd�l�\~}2;İ�諸��`��olX��M���K|�8������I�����U%��O���[-nm�/|Ȭ��n����n}ح���;ݾP�m,�]��[8���,�붪��m��O�V�ެ=2+^���Ui���D"�ʣ���k*�&�U"3^�c�OJ�G�-z������T�������C8�����Tk3��A�띣\�Қ�s���
֬
�y��,���G�`���}�!to����	��*�w�ۈKs��N��J�m'�x7�#^{4���S��;w������K��g	��y��L��
��0���}��I�M�I\m��6��~*X�/֋���/T8f�]k�t� ��Q10��֟I�׫�0
������mL��:��u������Z��C��\����78��8�I%����x�VRi�G!ER�:�`��%ذ�OG?ڔ�
4!�-���8�ש�|�7$�E|ǎn��n�<�P!=S�i�!˙��߉��ܚx��D\DHK����VK)��\�O�9�y�4��/�FŖљ��r�G��`9^J?:Wu!9?
�<�1�� w\<�Ҁ#K*U�_t!�E6+6�&Ĩ|J-�Xw�|��m�u%���*j,��*J�NOaHyh�a�v~��ĸ|Hj�}���LW�`@Il�:�,�t�PqhB&|�jq����*��U���腌���U����j�4d��^;^���F��L�7�<d��}?��&4�bB�֖�N��#1N7��$�e�m�#�4G�i��53j7��i���	&^I���^�0 Л_��Ŕ�e%�xa��閭�
2��j��p�et�̒�J�:�ű��Z��c��0��	3�XCJ�Fr��;�f8}��x��W3�Ft/8�J9B����8h��_�@
���4mm�w6�n8�闖�<�<r'w�X�|��j,�/5ik��FC�����C4f �,{����𽍑0��Ҙ#?�,�/@���a�p ����s������]���g�� �'#��K�/�.�vGaP�p����3��Yº�qL��F��g�)	��	����o[������Dd^�B�!����;�_	�ۦs��E�o�+����ڃ�e�iXk��i� x��Q�	X-`�	��
+��3vw8m�̡L�S����uK�_�Dg4�=�;��W������QY�6��v��Wn��f�RJ�f���R��(�z���#u�y�6��;�B��Ur��~*��[��epV/yH,��'�rO�܍Z�.��&�I��*�M�ɮ� ���v>�'���-�w"a��L\nʴE�F� �〭[��3��z�hQC�� ���v!j�T�R
�^��?�~ʣ��V��F;e
�'�u�J�n�ۻa�\&��mW.���EЗ�����G���uQ):���(W� �;���._Օ~�x�M}�1���������7����&��
+Y�/衅�]?ܬn>�;^�q\5E���Z�R�N���Mb-�>ׁ��X<f_�W�>>}�66'���y*�F�ki��nj#����偈�J�'�D�;_��0��������߮6�)�??t�g_�]Ȁ���� �pb�'S�Hq���������CI-�kH[VS���ao(@�Os�R�1�1A��%\{�㹢�.�jr%t� �ce�!b6&q��k��m!�Pd9��TO�H�%��Yt�d����n;�QMf:�)"�G�41c��fQ\�c��ag�iiO���p@��5,s�|���j�U�{5k��ݣ,�x�5V糦��hh������iL�'A�b�|�iz���fU:|V��ȡ sj�)ܠ��c���*�ϼv�.ӧc��Zm>ӗYKC7��T��#�-S�uZ��ZN2-_�RD����zE�j��)�t�(u��, ��B�	4�:�^T���L�8�~'Sׄ�y\�ª;G$z����nsi��߯8v����'P�i���Z�}S��Ǡd���p�\����q�)��w�V aL.	6xN�R��m�\I�Ҏ��c�F�g�Lm�]�����(�R��,uٞv˽b[����4&lzx;�$��6�~������@�al�cS
������f��C&!]�sV��IbN0��J����9���(�y�a#�]P���o����X�Uj�O���?��������>5��F������,��������<��"t����m�ßXҏ� :uL���O��(��r��)�x��� � =�qJ'p�Q��pc	>��.�����0ȔC�q�+a�?��Io�������;��4ȳ�/er�� +��h�Hɠ�����ͳ�k:Jnz����=m��PsS{z�֐�K���a_����%��� ��
���+`F+����pfZSNU�T��u�Ɣtc/N{�\���9C��3��.]��U�ܽl_C�1��y��gC<���yq�f��z4o>ݤ4#�I��n�"Y��/g���/���/���%�r��U˥6��"nl��,A�2U�|Ip�d�-8uX�S|�,2�L��7Z�2T֔�����e���ɑ���:p;�����\.?�50����|c0�ߌ6>�oѓ�[���^@�o�d)���vK�W�V�t�H|Zi)@�G^v�s׬�H��C��u�X��x/sڿ�t��¬���)�}����L2�ϝ�F�R~] �z�A,0A�c%����A37=ϥ�=����Ō�p��s��^�M@��՞CVl��(=��$�t5�X�ů*��~��-t2�*ݨe�"�1���#�pK�u����(u�9ٙ���~`��Y����}ΰ��5>�*���	e�\�`�{
n������%�F���ȊP��.�Q,f+��w:���2��c��Q�6��ܶ�]����J
b��Z].ٰ����²�>F��<p�-0�Ŏ����*�F�$b�]6�upq�O�Q��E#�8�^u��#�>8���A��Y�L����q ������ShZ�*)�`�ѓ��R�D�<�q�f��ý?@�;p	ύ7$;��s�mW�� L��^H(�>�w B|�3�����?��3CԢ��\X{�6ηS�a�1���im3)j?�p�F>��Y�2T����p(���+�&�?/����VW�r�c�uS�_���Q��K����&R���6�R}����������O�<�q�� â���뢡t6B�<<��R�5ݼ����3���B���x�uk��qC���8&f�����KK R=�5����.iQ�=��EU������m)��R��v�	�MCf�SUMr"G��`I%��]jׁXTlD%\��"��U��Ɋ q(�w2a��m�hnY��L�Z	��Sg���  �� d�um���!\�ڪQ:�'�y��6���a����8Y�:+%h�'�6����,7=׈���<��� S<cN�cJQY�~u����?��g��m�WTi��S�<�w�����Q��{'����H��%|��_�1�¿�=e��QY�WE�bG�����v�%�ZnXy*�C���������z�AH���\p��7�a(�r��ܘ��u�E�]`�a�I�HKb_��DL�͆h �d�Ĥ�c~ag^���4rd?D�?UU#���K���q�T��6��j^��\�9�*��"U��ɢT��"�����a���n�����^�}ο����x�W�C-������j
���I����
Ӧ�MK�	�_��.D����Dӽ��@���F»�t)Jy@�̐���i�kL�-�XT�a+)>����H���������H �)�l?8�l�P���;Vgzi��/E�{M����n� "+=�j�AJ[���DW�oװ�Ne��]KЭ�-܀���^C�w�AF���k����F��&��"�9�T��/zϵ�/��1�Oٍ�J1���7M��r��1��,��ómw����4B!�,s�v	Z+����������QZ�orA�s��޷3�_���Y�1�V�VBKdV,����M~Y����'Rq�׏�Y?A~k_)U`�\�co��\ ڽg�M]�f�0�]_d0T�J�悏y5|%2���;�͛�TJ.:"Н錥x����M�d��l�׋ntJ���68��6:���4G��s�kHI$��n�bJ:�+F���<�+0>�; +�E�S���&���"�5�W|@`������p���(0�ɪ峸��MVz�a3�yb�Y9wp�&�W���Ey�U�59Td DM�L�A�&� ���yDJ����3�ޤO5��ӗ�=�fг|�ѥZ��~��ʹcۗo1g��T���O��zx��5�{>>r{B0���9�f��}���=�O�@U�W��N�<N8E��Y��zω��H�BSI�����̞�)��S�{V��y"��÷?qLNx+���9�ʁjN�OyrS��;�� 4���E�0� ��¹dV@�?LS�Ij����P��9'�ٰ�'�2l�f����3<��Ys�(
�I�⭕��E�#��*��\�9j�='l{�`3��5$���	����H)��qr�J�(W �Լ�� 0<����B��쎁���0Z���u>��G��tC�b���m�H��t��Xo��JM٩�ďS���$��ėmGt�[�G(����MU�R�U\݄�¾P�6�`�8�	����daS�*-XK����d���!���@�O��QM��5f㓞���.�t�)�qzZ���P�e��AѪ��(ӨD+목7$7�x���t �܏�lřr�{=��m\s�6�y�{w.@s77����92H)�P�]f�Ԣ�N�%
�;��&م�?�L��nÃ�N�:�*=�H�-U4��;��	������ߡ�c]6���`�C$Λe���Ւ�JS!�g������l�9U!�!2�ԛ4��R���w*\�=�e�9�.���	��5&΅�(������D(p-��(��+�LUfK�5A�~�`��@�n�z�,o�F���/"�2��FmdZ�UY�:"��D�[��[ho"X7B�~2V�T���d>tw/g�t/.m�^���ߤݫ$��W��'�#1���4�I鑙�5tu��q�% S�T�e���reU�L��7�$&��L ��?yC���;���?MaQ�-oP�L�D��w�ѯ%�+z�s��8��}�B��@Qw���Ƽ���p3�w����3M���.�;���(�'�i���;R�z�dN��{��sc��g�6Z�%���W<g<�Kh,�]b0���F��jy��}��i�,�j�J4�8pٹ�
����Qzq�'���1p��W�"���	X�m�'��C�����J7$��rjek�<�i�O��h��s���o����c�����5��2%��0ԥN	/�#�#��C�ᬰ�+zU��^N�=y���-+� ��tL�QiOpnj]�'|w���3� 퉋�y�~�M`m����"�]�y��v#����۞�9�{���O%�EƸo�f=E�w��J Ƭmt�n��.G��ķ���;N�~}�����n�n��*]����Ws��)��G�Ց澈�� ����Y�=�5?W�	��騩`�rH��:V�Ύ󱘒�Q�"|�9�5t��|@���{^Z(��D���Հ^k���y���+�5Yn����`�`��d�G��܄I����[����L&�z$1�q����᫆��1�
�5Q���;��5��H��yv7X� �l���Y�C�2ɱ���J���Q$v�C0�x�Z�����=���2M��%�Far�@�p�Ngl�x����@k�U�|Z2���j��ύT
��>t��p`����c��z����%[�`��_�]܆���XL������t�yV�|��#��wCT���B�]WZ ��������lz	޷2��f;d��}��g��ѫߢ�ʮJxA��@]�,@�U6�R<RI;u��ҭ���_)��,��6�ۗ��9VJZ.o��9`υi���T��C�fΐ���N)�Ŏ�e2��Y�^�n�{ 7�,_��D�~j�&v]і��)�I����|Z���E`z��8Eb����D����3@O"��I��%ЯI2�ȱg����@mg"�1?�a�f��o5'%(��'�W�'A�����7WfC�����@"��!���ƪi�ly3�^���l���J��Y/�#;	�6����Sp�
�eAK�ݚ?a�d��*e�xZ)�"����ݙ�Ԋ2���w�s���`��3�m�<0��`�B6i�ˍm�7<~�0��{)W{�8�[i�X7�&����N��Q�_RP�?|`I�A�
����?vƙſ �^� �e�oH�5g�t�.)��>�a�%�QV�r==��ư7a�ߜ���7-��x�n��M�C���ќ��bfNf�@7�����0ƪ��׸�y	�X8h{DE����U�a^�?����n���~)B��Rnc��|�VTQ7,L@\�B�;�n���Qې�~���0�k�Mi*�cq랿���B�֥3���:�Y�?�=f���ڟ��sV8R�Ǝ`�M`��H���5+HjWCl>��Wߧ1r������1�6a�[�i����V��G�%Bw�Ƞ�S��@NX.
�����&G��m^$��U��7:8�zc�`'���[��߼c�1"o��z���fy:$vX��iD$
���B�$;�<���*n��P�����B��RK�&�!�����k�x{P��j4?��2FWcSp�0]���C�L�����*�l��+��JdbӚ$Sa�`$>�T׎�;TE2�g��oW#T�M��5Th��Q[
�N�u������a/x�p*����g)'�@;��� ?���(el�-K;�*1a-��S\F�#�H���6��G��I[��^�óS<&$�@���o�_�=6x�HX1�nV�t.����1=��M_��B����7�-�}N���~��GN_����T�=Mѷ�,sy��cwAQ�g�"պ�G1�F�5�����J`�SH9Rڷ��TB��k�h�8�n;� �t�4a��[�FP��U����cݼ1J�P�1���=�]=��>����ˊ�{���<G��PT�db+9�p}���8�L�x�y�9��<���҇�n/�O|V��Ι���>U�Zf��1)M�����*(G�J��mk��?��g�obF��l��4Y��`k�,V!����c���T�c�� C�s�>��{~�;�m�w��+B?}�����P�7��n����5܁0�a#�vx���[l|[��c�ek�d���̘,d��|�ނƉN.����`�?��ASb����5��o]�mx׎a�+�<��i˽Ut_1�a
W�~���c/�C��W���y]�v�s��xO���]�Л{�'��s ~�t�1�K=��.Ρ�+B	"��j�;�S�īG_M�nN!vU��>
9�43��LL����/L~'��g��X���h���?�V8y�;��)0�9�0��!6��qr���
T�Wo+�+R�6$�����0�e-[�	.�3�*kǳ�c���O���A�9�XK�d`���3֢�9w�^����Vj� �	>mvK�J�^:�i���/���o(�XTc�f~;��ջC�۱E����q#�����p��`���;;"��z�^L����o�ܒ<yQ�k4v�'V�w>|�*�}hS�ڱ+Ӧ�>���J��߷�&zs{	�����X�O���o��pP	���aYL9�x*��G�'ZI2��nr.{�Gh�2�Z��ʧb� �}M,��>k�A$J�N�ȒB�gt@���xx�_��v e`k?�$��$�@� ��@"�C��wN�q�x�m�d[����U\�|��aGt7�u�D�֗���^r�w�)�rY�d����vq53�7��T�7���-eWK����s�]L����d
��\�`��)ͻ�3IO#7�T N�_�Y�[dZ�������\��o,�d�L\uԺ���}�� ojf炡�������X���[h�Lِ �B\ ��/[�6��eYh��<�<�H �)�(����/�V�W8��V��ۓ����6�	c$eb���O��*P�L"7iCR��N�ч�+��}"4�_D�W>��*!I�e���P�M'�)i�/jt���Q_q7�)
=�I%��g�܄"3�M�DF��sR~N�طG���x*�7@0���D�洘����eٳ��e�ߵ�ՇЍ*�(�L����Ьԙv����ƺV�{,)��Yh��g�W��'�ib�,����,4DL I�AXT�F4{/_L��t,r�>(��q��Y��V<��XO��P�eE5V�H>�A�ȣ����� ط�N��T�B﫡�L�?��V�8�g��@��G�6����T)�(�Z�^�z�r H�9V$a��W�i����t�c�T"�^j��z��F���2"R��S��^wM���9Â3�
 ˦���,�X%�C5V$]�M��Q �4s}���ʊpkʿ��OsD�m����.T��Z��C9K����&���ƺO�a��rQ�W�=�-���w����]����i$�v�C;�P�3F�[�~G!�7/A�I}~�� n$���%2��Xi�q�	�,"�mI):Q'ݞޘ�J�;ɻ ��×�q��[s��Duds��5�<�N?/p-hhl4>�?�!�S��OSi�]=D��� >��& �"��Tt��f�~7z��a���@�5WБиp�|w�G�)�'�,�p^�拰UE�sJ�Z�.h����\�O��K��u�M[Ք]�+��{�=�[3|�=ˈ��Wc�SM$sY��L��%�"�5Ǘn��]ݯ�6�v,Ձ"����f�p�C!��g%�X~Q�#��ϊ9� *�d��=�<����%۝��-���y��2�7�&Y��oN�����s�y���z�2W5�u,{��d��йI��=qG�O�$(o����=[�4�:���N����j&����;{��+����ӇNХ����ݔ��I��]�O�ƀ����r;�u㠲1�=f��k�M�k}�|��&)B�ÊQ)HX�Ø{;�	RCb겥L<���>'"U:����2I#�͟�!&�^�d�`(��dC�S��+�bf_M�n���Q;-�����>z""4ʑ���	��� ��.�x	���<<mv��'��m� n#�#_6�`�y�&�	*������K0K��ǲ��M�U�G�VYC��(�~��(ҁIj_���o"P�$��Vn�L���R�q��)%�qo�����&�Y�����(�O^�e_���}Q�c�P��yT~>@���|��(�*W
{ti�û��m�s�*��S>F��ş�
�����g���dQ�1����)��L�4Ы�0LOu�Y��s�C��*�+7r����]�BB��A�Đ.�&�r��2h�u%��q�{���Y/Z=���t�B)jn�1�;7Y2��Nf��hA�x���ܤ����_������n��M���0����m��O���x�j��8�'h"����9�ӷ����j�֚���f#�x�R��������ַ���6P���K�qY-D�ioL�x�� 1xrb�;bx����7�J����m�:r{5T�z��d;�B���ٍ3;��� 5H�f�f�� ���y��
fX�^/��)���aU�F�|�I���.��xr�r
� ?G�^$.D�,:9��y�A���C���S۠�nu CN�%�4�6���1�й�]d��j�HQj��<xW���˙V3p�t����]l|�eGq���-)<SQE����~����Cj�@06',�P�֘�̚h��%S�,T�����޹9F��B^�]�Jj<�'Y?���Tb62%��@� ��WT�]\N�P�%TޏB��;V$�Ylݪ�d�PMW�5m"	E,��'�@�|X�����dSH����|3�����:��k��\��.�E�u�����$0f�Φ��� ��#$M�."�?��/��'��F�Q��������F�ء����Tv��>FA���/J�艥N���Nc9O�.�u�E���'V!im��
Ÿ�ۀ�:?�
����Q�q���Rh�C:\��(F^V��$s�j4�O�ߜb����\6I���5f�F^os��L(�3Y�o�ټ�4E{��0Lƪ��2�*�ri�8��B�J�Q	'�"U�<�GM)}gN�go:��풜�-��Py�+�%Ӎ�8x���4O��Jf�a�Voc�5H��uG�=2X��E���ݽ�}�OG���wfL)��@*���W��¿m|	2�YJ0#��
�։.�X���+&E5 (3��)���p���¡�ڮ�.����dq�� �d�C�8�ft-u�7)��������9`�q��3��yL���Jw*d�zŠ;�����Z-�?��4[�N��	,&�Ӽ/�E6+��`�u���;�H��+Z�(Z/AD�3��)r��.8���B
��ǌ5q1;2*��Hй���N)a>�܈�O1�A�^�<�+��y�t����ZU���1���#y��4��
�V�ރ��ʡ*$��_��;�1�Z�^4�Ko�4�-�>+�{x��k�v�UA8(݌��Dˡ�ԏ�xP0�4�'���t��x��CN<�;;9����hA�Z�7FZ�Ɔ�L
�;�W�fw�Tvh�)�{��U��k(?�P�,H&�r����=�]���_�uu����t��Vՙ&h��3}d4�'n��HE�u4�=�O|���cͪ&ey�f)�j5��v?s�2�0��B0��b-���?7A�E�5E�긬9�#z���xpyW� ��I�4�2�l(/|�5�gA�2i&M�k[�����o�N{
�XX"+�t�+�]g#�֨Bm�?4�3F�S���@���0/��<�w���]$���д@��z%L\'�h-��jgZ��}{/�<6m8�e�@�!:�M�����w�R�ba2Ğ�rU��b�(���M3`OH:�ӫ}�҂3�����Ţ<�q��!��l!��2�Ѫ�Y��k"p�ƛ��m(;�^c�V�	���ܫ��4wP)�D���^W$уD�蛅C�U$I��$�uA�چ̠�cJTgRT�`٭�6��6?D=��qN��KП���Z�v�Xj�=�-�lj;~� ��ό�#���L�5��`Cbk>UA�K£V��ƀw(Q��j[�Y2�/L��HU}m�K�b��`H}��ri&�4 ���0�Y�e�%�Wx�qc�1����=+��G�agٴc}/�<\�\Ϻ<��L��_���o��t��ZG�k�c�>J�/�J�HE{s��n�gW�+
@%Y\ݴ*�Uۇ*^84Sqq�~#,��aҸ�:�}V�A§�4�ZN���>=�4W9#l��y �O�|GH=��ƭh�����)��~R]����|T��V�S�{`a؜�y����s¼(y�X2N�>�P9ۿ\n�<��O��ÐE�k���[lTAz��*i�U4����
�]���_&6���ri	E�5���ҧ��щY̰�գ{�>-�^n+��#��IYq�����R�$��"��C������n&�ik��8�a���z���D����{�[QR��_��*�a�*;�����+p/��{Y��yӟRH�ô���"v���>����ͻ�K�~hx���?�A2_���eko\�/��6X��& �q��.�� ֽ�� �VU�fS���Tl��=�2�X�D�3����qD,��X�j�Q��"Ū�)��oC֒s�;V�_엔��$���<o�����=����_8!���Oipި9%�eT�:��B}b	?���?֛�}]�º�}�J�((��-��`�����;��rd�Z\�JC�䔾�# '�Ae�pS5;!�C1'Qa2�_�lk{�u@[Ke��)�Ґ�/#�Wɩ�?�*�j��k�v�V´%�_n����̤��$OT�%�J%��;sM���Iui<�q���~�7�q;�6��'���]$�X�(]��Ř����!�ϼh2��v�|n�u��K\H�J,fC�]$6��J�UWT�Er�z���G���C
y�/���]t�$����l{��5o}e��9;w���eo�q��f�1`��,���;�}�b��U�	 �6��m��2�p8����L�����Ԥ�Sǔ;���8�ƙ��ǲ�Ї�� �\qY{hjF�X��$k�z�9f"�O��>���R;�H7E-R\�� ���^(���W�w]	�e�g�).�J�f��Y���w�G��	=f|{����y�����J���a��Bt�HW8o竘�+�T@Af6����r�sR(,��U��UmE�wM��(.�c�bɫ��N��ᜫ�L#�^9�޻������a~­�.-̛c9ESEY%F�2�f�r�v�ՠ&������|=�J+�z=����C�R;]�x_F��d��,�� �����3�ȋF^�&h	A.�:S������^z�%f��J$�0���3�5)j�JQ�&H��˃\4ӜR����*S��-0/Ϲ<:����f6K��p�
���_��-������nJ�s�l����+<H��z�PF���L���c^��?�|�`gT���b��wW'R?o/:�W��� $Y�
upn6ʑ?0�KR-HH�4�X�vj3�
I�+p�j��u)�3oa&}^̛a�3��(�/�1�3:�Lи��um�����Ȩ&b"�?�,�	�Cf�f�*�����\���H��p|د{����ʢv�F3I�V�E�Aޘ�����M��I��ѡS���Sǃ�@�m��9+x �S���4�1��&И�с�2Q[��`��j(�Z�R�K����N��u�G�Ii���jE��p�g�D�|��\[��Ev�zOD*�'L4���i�ŚiA��v�3�)Ѩ+1���]�q�6_���g�$oj�~.4	ۚ Yq����7��U��@��L`�~#��l|v4%c��|���MM�ȴn����ލ�?�F��9Ӹٍ�b��	݇Ȃ�k#3?�"�{����Rȍ.P��n��@@�� 2�y���m�7d��{��TVYZ���7�D��n�x����T)6+]���뇉��Ⱦ�j�xq� {;M�B*/zeԶ�i�L��d`ٛ�B� �K��ߦN���zm��C4|PխB�3O�	���BЀ�������!��w���Tnj�����}dwS B�&ꛒc~��_.1�WbV�y�L>Wd�[յ�]�%K]�7V��Q �Ӣ���ΠeճG$�u4|t.��W`{ݿ������`eU�2AY� %g*YO���!�}i1�Yı��X���7n�ȑ췚1=|�ol���[Wy㦮l�CE<�h��J�ғ����V��� aӔ-�0��Q��,�䯈��n�'A�,�LJ�6I�6�|Itzza(,�Xl�i\Ǽ�=��Օ��&��q�f��^ȃ{�ڋ�)�ڎ��,>k���\���'��Q+F
i��
�Mŕd�������;UP���ҡ�#�z�KȦ��a/ ��ri� Խ�G����盗�OF��Z0+t}*">B3�ĺ�=��,�I"'S�tw*n���$��MD���S�4gi>s+M��.�Gu1RM�ܼj���e;@b�\�.��cھ�S�0_��/@���Pe~9o������o�p�N�XUr�-�I"Bn6-7+C��~��%�Q@�h%��U��u˛}b4�6!���n���ș$��\ ��{a5h�NqS10M��Z�3���q��d�}��n,y�Hx>�<t"�>Ŋ�ݮ;��w΍fG/.~�k��ŕ�H}��2J�� γVM45�(�ڌR�R�8��LR5٠y��r7h�Ն��#�j/�
��!��YF�B���̈�	4R5@Rc�����wU�1zϻBN��A���ϨD"�ܑH�A�����H����kF8J�U�(�)���J���l������X��'D��%*z�l�x��a$�6�Z��V7+��TV<I`�+;Ͳs���u`��1��������%t�&���^&?�d�w_����A��#>Mu��֙���#���µ����H�j�|�8q{{�_{{s72�1�:����[SH�|���hګ=��Nz�t}"�EE��Q�m���ɝr��voH�A�Q�*}~	G���J�vh�s_�	�P��Y�i�������aA���)ҪU�� �ِ�� ^�EJޯF3`Mab��Ib��bsd�*x0b�s)��\":�Ԕud�gثQ�Ա�p�$|�N3���h?��������m�:�;�qg�ᗰB���dd;t7tW�V�}~{��Q\ѩ��"��I�b��nH-^�Zֈo�E�O*��#x���z$S��he0��b�\3p܏�s-_�$�^M����9�9��cY�E�\���L[��7m�yzF�5�ж�Ps���6}�-��ѧb�Nx�$b5űd�42�.��Y��N��,��E��Tx��aa�-ܜ�o�T�jn�\?갭õ�O��L��Ҫ��"v^ļ�p~<+�e������c��k��]$�B)�2�2hHJ;���5�J)�`�s9��~�#~��P�}?Ԛ��4��M+�	/�c^��j_��d�j$�;4�g�D��h��@�>f����x ��5�&���� �
t�TI�6*��(���W�?�Z�k1����bL,������)8ӂ�ŶA��2T��Ձ��݉���}{S r^鳧�|uH�̰���ߪY�ñ��zs����iK����f�sG��A��k�#����(\���7�s���s߳�����X$�4.z��]�.���C�&�b��;��En���嶬8ff���p�y��=�ܸ<����
"�������]=W5Z�{f�M6�ꍾ��+$A?��ƀ�t/�D�����疓�=�\rG3�:U���
cr��_�uҨ5�����e�q��i(g�;��^q{�&�E`X����.�}��(��D���������.@Z��Q|� ]��m��w!���O1Nf�����2u7YS����������$~����Kئ.{�>��� ���[;���T��V�Ux����� �2�t�]��۝�=�>9�I�1ǵQ\J��۵�(�>��~Z�W�<.�er���m��pl���MVW���	<@�%V��0{@���$�W��#���|����0���d�JMg�A;��*sUtx/��)����?[��E��(�5�ϳ��K�ېuo;+;��pȿ�-��b����PR-+S6����˂�_v��y�^s峁Ey]YJD�T&����ﲲ=��݊`��뜘��D��	8�a+!+6c����o~*����E�IJ0�9�E'��@Mhg�ڶ٢av��@1�GX��~Hv�A�Xڎs��l#Ha��zIr�C��a/��j�;��LMe�l2K�γҠ+:��y���I���"�Q8�a���r�X���Z�'�8�>�X��o�F�p�Q�(j������ҭ�����)�t��"����	I5�oG��R�f*��L�S]3�b޿��RC�`������9(}w"��L���j/O��VN�ֹn���5TSD��EDf"'S�_�������^l ��y@�5Ń��"N��@��U��pG�e:W��BC�?{EN����|�w��M���y���9���M�Ij�oq�u�������o�BZ�_���Ϝ��bv�
8e�70ƖyX/���D���vD	F�����.��F;E�᦬;�	������*1)�ww��	����\���y��(��H����@��&$S�g���t�[�/8����I���/{#�L!`b^,TG�A����S�/�=G�y�	���n��,��UO#��$������Y��o�8��#�#5�#����(W2LZ$��':�`�s����	�*0>x��x<�������p'�3gV��~?����@U0H��A�dʹ5�;�;т#͚J��H�j�����r�"'j�bH��Cn`�@俞�(��jQ�������eI��4*�r���Z�E	g$�ݩ�i%m�\
�j�B���I�o}B��m�M�\g,"�|��M�6�����)���gyy�^�����rL���s��[�:��R��U�H���_Y�D\� ��T�m������Y?�w��Vu	5�G4r�����4����`���l�}�{ �n�W3��M�Zy�k�a��D���m#�!��	M��²�d8�敦��i24���D[H��q�.�:���2�0W{�������wJx1f��lZ]^���!�'WQ�����r姉Z~��vd`���EG�4�,��X�Y��B�t#���8��瀁W�,5�&�J�a1������a�������nh�h���?���pہC����]m�2p�-��*��$\�]�B@�-/ �RxP��(1��3,��5p,1>1RK�����m�O���Ǹ��-ո��W�ʊ寗\Q��z� ��pXെ����
ܠs��+A�_�U��XS�hjR��w}�Xf��4-"@���]��P��-���E�+SK���`ږc�H��8�΁�V]�ٟŧוB�lqFlä����br�<�XD�c�OZD��ɺi�����{z��� 0´RQv���X���j�	O� �Z���w�y3oS6�hE9	�?��^���ڥ��̎4ƽ��7�r����MM�hE��h�z�p�x㸻��7N�����7Sڗb��֧Kz6i�טC1!4��;c�
E�#}o|���Ĝ����s�I�;���	�<�{��ޅ�fQNBX-�	//�� =�T�e�]��W�v���uP�\��\�..��o�y�j[IB*�|�������E�w�`r�FbX��}? ǿ ����Tȣ�Y��>v(-�����Ly~����a�`@q�o�@�֟7r�/��
6����0diB`=\
�K����� 7.����ࡤ�g0a[���T˨5b��j㉯����V	��Bb�i0�`�E��AY(۷ç��ꚝ�YMӓ�y���ֿW8����G���> ���_���,Iş��!~�4���N�����rq��Z�m�lA�&��䗷�x�&���Ka,�Jʖa�<�𖧣�'r��1y�r��\������=[�R�e�*[w�drω]�i���
)h��_�=M�n7 �Ǹ�����<�`����-88�X��F�Ap����9�57h1V��� �A���|�&�T,���� �д;K:�v'Dmi�;ޟ	׏:��ps��?���L� �����9�K��CD��(��%��QM�YᄷB���;͹����?r���LS$�^Y�zTN!��u���5OpѴFmf���b�еQbNLR�Z4�`JE��%N�X��#Jf:��cY�d��Y>�~�/E�M����R�MAg1 ��J	��p�@U����|
��6���.k���7#G�b��q�|)�J�>���v�SY���w�E���0��٥B���G��;����R��t���&�'"{2h8%K����S�ב2f��M_Q2�f,���g��N3ڃv��1����j,���B��I\��z��_l��-e2�F ��Ѱ�V��硏̣�Z��8÷>Ѧ(:P�	9(�s� �TsG�/QБY�"n�\�*P�%U�H:@>�|���Q�c{l�;��;�sҺy|.�a�DK��a���?ŋ��0y�Y���ߞܚ[�G�@.��it���	4�{�&��Y�oyd�J2���k����a��U���zE���G[�ޛ���`���邮� 1s	_�ֿ�IB��u�Q����9��
Z'���Âҙ�5��bU�1�!�	��U�A}M(��HS�����;~ԃ�YҹI$����j��܂�9��B�X���~]��88[������m;�`��`�E�­��bd�MZu�JY�#9=K\%7/Ԉ�/�`yl?<yy�}�K��x4��9ò]㇣x�C�S8�-Ż7x�O�ѵ!3������a 6\JB�-Ѽ�ޖ�-��*����c*%���ތ%�Z6f���h�_�[��q��dޡi���7���;�fbk��tϽ8m�_'�P�oVh�W�{Lx?��4j�1+Ҕ�s�r,Hd׃���YqK�֫��@|e����-���Ǆ)��E�jJ4!���\�bT}�x�ۣ!B�d��핥F���oK޾���r ���(�*n{�OF�*�ؒ�6�[�W�luN��t]Zl1ԛ������Ϗ�`��\�^Q���f�z��Fl��L���<�|��2�퓨P�x)��1�sTA7k�	L�	Xd��
�`�6^����)\	{#ta�]��S4�F6�&%���S=
��.�A�����RH
�˚{³�[ժ֐�0�;5���M��|F���ރ�I��^z����.Ɇ�gÜ�HO�I������ږL��}�n�	A"�B��m��}\!���E�xm!�_z�A� �$b�8{��c�_Ö�������e���?+#��9��y^�2�#gfF�C��Ǖ[;h2�a�v�ǥg���u�,�z�LÄ:3�^
�Zz �Ң�wO�ԑa`���I�>p�.�=j,ǭ.̹�`����E`��ҷh䪨����4]�EqaT��ԁ���2c���"5�*G�O��x��'��ů	�Пi��즕3= ?�)�Lf������f6��d��W��ca ;Bv�����}��Bo��n%P�#��u��N��gٶ��/��
�H�?B0�Y�*r�L;��ݖ]3�.c�h��}E�K�pKq��@u��;<�`����3x�VY��St\��# PZ����0yeϪY�J��)[$��$U6�T�M�����NI�T�Ш���'̛Յ��戚�Z�׆{�����Eļ��&vy�Jy]Ht�S0�XuW�
�?'x��9q@��RT6�hFMG,�pMu!�"�t>
l�Q�S�"��+k�;��C���)r~9/������G=U5|y
��0a�٢�tpY %�hw�/���JRc][.���w�9��Πi�s�NA|4�������ڻ_�V�&]�Β��������g���1�к��n*�H x�P:�(�����a3(+��t=_E��0*~�k�ց�w���?���Є~6��9���]��qMo�ۢ�E������欬ᮿ$�ՕC�t�,i�s�jc�pl&9X��p�]��_�T�A�VH��$8Ǻ�,��]��;��#��a��m���S�m�3s�e�2~DG���U���|�Q�@F{���f-��]��qQ~�rWH��^d���x1���{V�4��Hjǈ������#�ovKTrc*�u(#�5�e���xc���a����]�̪���9��5">Wm���^V���z��q�YZ���ӑ}"f��d�
�Џ����`���2ō����*�Wc�:�-�оm��d���COΤq��L������ţ�,���
�I�2��`��h�X�c֖aw��.��+�o#ȩP)|�(%c�5p�5L%� ^�.{�w�`H��ӡ��BG��q�Q������6�殄+�*rc-���n��D����T�8�_#/2m�#�z�AQԻ�l�?�ouRI��v�TG�Y8����kw��]�I�B�ꇿM���>�Im�R��k�ca��ZuP@	�����z�s��e��jB���M��� +x$5�)Y���t	j�IwB���gN�1)6}�CkM;y��QHd�2�/NﬦD�cE}0DI�������-���kh�T�=�m:�/e���	e���i��;Y��D�`��"���v8��c��~��1���]�(�?�����{x��u顲OjM{�ޒ��ȖS�q�
hO)�X��CL�����5�2(=�)i~�G�%�[�k>b2q��F�r����+3�V$3�<��w�q�*F���s�搫�4�Qib�$FG���j;�`��}��r��^�B$��A
�����禐��33 óJ�g%��Y���Ԁ��6������{�?��$�"�xc^/����o[�\�{wH�xtCKG�VH
�nR����@�Z(a� �q�y؅ר�S]��$S}���D!�~��UbIޭ��
��H�ZB-3���̚�'t�?53��N_Z(��o���������k��{>���z���៵���]��3ጜ�YlH{���ݛ�3�\۫�3�*pB�'?���{���lNc���� ^�SB
b���^��2W��'�J<4�,���Un���}Z��.�N�G9���/�J|�n�� Q��=Br��a#ɖ)+\-�4?���V�����!D�9T0�#X�+�f�;�����>��+��>�tn(�X=7�=u�R�¹n���ʸ���:�"3;��:H�n�P%<)k.���,r���}�J�m@@h~��,K2w:�
�RҲigЬ��p���hB��Z/ Z���Țj7�h�z�w�0��'�#��S��R{�ė��.�ݖ-�\����z�R I�P0�����{��;��j^>
lWM&#�Z�M�>���y`�C�?9ܖj��25�0�J�;��������5���vc�-�7q��w��:�@+l�5�`0�졅���;���Z2�#�Ю�V!�C�_f��I���0��hg	>ՠq3jl�#�>L�E�Y�o
���ww
4�[,tf�0վnԻ(aęv/�ag;����D���ɿc~4��i>u��RYB�	�~�4��c��R̰[�����-���B����%*[�F�o�s��/�j�N�g��s M��0q��M�|���<�Pپf�n1�ɉ,�֖�/�S!�Þ�d����m_jm�k�_M�����|�����{ �%����2	$=U�L�qs��f,��H�%U�U���3 �LWO���l�k�bZD���� F����ʩZm���l���Չ[1/3#�2R6�h	�ntOc��E]������_���O��v�	g��á��%��"����6��I7G�=iOk�p����so1q���fOޥ�I��ƶ~����Fʐ��d@3�%d@Q�060�}&:s�
�@kE�N�5�
d�����k��TH9 o6}-a�MYgؙ9�[r��H���K�74^�k)�	~���;�H����M�}��w�45 ~(;��?�o̹�����R�P��s�)~�9��W��`\3I+�Sه��~��v8f2����0"�p� �

S�-�H��{Ҿ�sׄ٘��'�>%B]YԪk&��(P&P|��{JgDs�@�	FͺO�}Jĵy҅���&�������5��i&)B�M]��Z�7|}�ne��9����,k�Y��P�i��?���Ɯp:�Ck-�dH��c L�=s�[8�zV�u��p��%,:��p�u�V��ޖ���˪hKfB�g_��/��C��9H���`����b�0 �r�"�}fJ��K��ß9�����R���h���?�E�*��I�a-~7�ܷ�o��6��e��A ����j�l�w��d�X?+8�"J�Y�J�4OcL��r!�7!LYLX�md�ޓ��My̯���Ki����dA3�E
�<��E;��T�0���k��Y<�0A����.��C�&Ϊ��_o��f[ÊP8Dϥ��ھ�P@O\�?��������e7PRy�rq�ʹ=��ob�B��Ep]��Lt	bD�*p:�ޣ b��ģ�����ܱ�P������`�ȱ�d-6*��T/����h�����ԭ�y�V���N��1o��й���휸9�+L�z�_��]q�w,��-������}H|�8���ja �<2�#��$�k\	IZZ��s}��]�|=���[�)���#ef�~�y����H#����B
]���%|m��~Z�������������D�����4�}{���#pX�`�ݳB����N��a*�]�vW��ӣ�p�����G9�z�Q�Hxjp�O�;���Ô 5<����0�ZH��.R���
U�rЇ�מl"ۆ�b<��Pյ�U������6� ��\EA���9�CKA�������rѿ1�������,�_�r�o4�t��F�+��_=Jصa���"�.4�g9l��P��G/O�j�Ǽ� �ԞpC�{V�G�Ҝ�t������!lh��烪J��;?=��j+ݱ�2���������v�C�n�5 �.���>��,E��A;��0���d��l_�^������Wb[L[t��{�3���}���,�Y)Y*�ծM�����q����.���1�˥.���_N�r���¯��8�Oˆ��Bh.Q���	�b���ۙ�爉
3X���@Q"0���L��&��G��,>�<��蓼�e��`�o��ǌc=�,�����|v����U�}1]�cXzT�פB!�����[����&p�8e��yS��/�j�Z��4	��u�䜜�g�Z{<�/Y�y8�Ş�8�9/$���"�	�$��o��u�����x�*����O'�4>�G.���!��w+�!�М)�M�'�ˏVvX�!$P�	��!幮�Ҟ�����@A�f5�h�>g�����ڠQ�\Ӹ�s�y��-��l�F���w�V0�Q}�����E�T\Q���a{79�eտ�܂�F��B�3�����睛�� Գ��l�p�p�rAIS��g�#��Z{��g�֧�+�a�0᫚s��:Gya�5����Pq���*�D�"6	��c���~Y7HA�
t���2��\C+��"��5�<C��a�����$Qg�$ឤ�Tϻ��'��A:A\�c���c@��������u����=!���K�6�w��%�o�H"���L�ԨHI&���K�ٛ�Ċ��s���b/t�/�M8����cذ�~!e�����I�6p��;q�73��"�-�el �	�v��Nf�?ۼ�e\���4���xT�cf�׭Q��K��d�%!�z(nԭԸ�K�'s.܅m�
&u��f]�_�����6�\x/�'�hO�1��IYƜԫ�)F��� ��*�D�7��ct���q|��'Q�j���4�ߘa�e�4!�t��:���g7�'��Q�B=�@��m�ړ��c&}��(9n;�j[6�4�q�\q��~����j�b�����F��'�}v�w���k)��&�u[(�0�����*4 �9�@O0���-�O�����:���䠡�K?J�z��z��͓�`���ؓa��_`U-{>+@�_IqR#F=c��#�ح\&�B랟2d��_�v��A֤����� ����Dð3?��Ex�6M;	v<����{����D�ס�7-LǙB��i��u�K"tB�_|�}�"�K	L���<�ք�Ol4�-[���01#ѿ�`�.�PX-����(z�G�W76�>7ɋ���b��$�_���v��r(z�ck���O_�����B7{�(�R�Ƥ1����x�J}��ג\���&d���bc�*��h��$�z���2ǲ/A�����$9Jihpƺxf�&���x���}�nHk-D�O����R/�T̒B}Y��a�
�d��E��T��+�j�p�'�Ѭ�gWv���Υ�ɴL���ܰr�9T��~�����͌�3��`2�� �~yѱ3�oQ'q.����1�X������PՎ;������a,w0����4W,����p�^�E�2C��"#ߓg��ʲ�)	�V�ڦ.Q��i���R��#m��*C�Z.8N�|��B䣝��� �ly�	O/��Ҟ���G��v\%1�hy�yc��I
.G�,,�)��2��h��&0�4�Q�W�P_C({+Vb����X�F"i���	6`-����+�a�,-�7�,QqЄ�F��T\���ڣKȄنG�-}?�n�H %*Tx�YX݀�m[�m�}�
?�Z^�ץ��jE?���^��±e��	�*�-�i�!�J��I�T���^�R�1����qm�@�6�xFU�}SO�@Q�|�ί�
)��"�ZV��}�-Eȼ����4^����
mP���Z�m&�<�Gъ
Pm�?��S2ST[�6HM�@�WBZ5�x<>�cd�$5���#�����#���P7i�i%',|��Pm6��r�5�n1��������^�ϺtE�k��Z�F��4Bq?�,.��0�fc�S&��MD�}��uj����,G^��UauE��6J�B�O�>3b#`��Ы>Q!���agWc��L���<���W:���XN�~�O��Mɝ����y������HX�<^a{!:�k�6��B�7�{���uCy�>Ph-j5�mq0�J��Ѷ�G2��C��{������]���[��{z�Tߧ�>w9�6m��c�VM��j��7ڼw]6����w�3������}��͒�el�Up�t��/��~�1i�x��t�!��s�V�|�Y�f�j[�����ڮ���	`�[�@U.�C=��M�	��yoOk�z�`�ǜǃQ�d����p��P�E��m�VU�aՉ�q7P�ǈT��0�7 C͑Z��g��}���c��&=Q�E�ޕ36V�'M��'/V����x\A�Ti��%��c�v��V��c��[�1�^�B=���9��q��_�A�ž�V�w9#��=��ez���|���/�ùEBp_=�F]k�x���s���1#.�m����/�C��Ԣ������,�ײ��;N�U�v#}�U�^��u�ғ�g2�J-�V��T�5��μ��˻\}r��ٻYɗþⒾ�Q>1��@n˻��r��-��D�?�O���:�v��o��%�d��hs��;`�V{��Ҿ�� ���ӼR��+��WF�/�޲C���X������k�v.I*^oE��ݤ�t(��ܝ��Dԩ�(�P�"}�%��`��X�'�1�+�?��^��0u�QL���-5���
�"��j��c�sS�*�JJK��S����84o���{����TB27oA5`g7�ɇ���@�>2*��l_9.��=qH�F~���;ʛ��	f|�x�8�bb��{���OuB�0�/s�s�꺯��1Dl�41
�����^��i9|��H�����eo�K�v����tŰ�����rQ��w�!|�Д1i�fp���pmi� �z6zM�ܳ��9��,�7[0m����T���f�
?�"�?Wlɝ����>S��g�i��^��ᥧ[��"
 o�p�I�J�T���`+���Nr�S~~@#�/H�d�����*(��s�7�͡7P��+T���o�|�T�L�	�YA��,���
�J���Y�"�P�S�!-t�P�Uԡ	�G�/L���8,�'o��P���Q�vjFRXI�� pVJ�}��s�^d��|An�#�m��cl$)��L���E��,�t#��hI��K��e;���6��7�z�}@���?0���P�g�L���I+_���	Cu�>���dˠ�1�9�sT��gԖg�	I�"Ƀ �l��k�:Z�fB�JYu1����z���:{`�3L�{��i�=��ݟg����*�;�WR�m��(ί�\U�+u�1�Nm��>���}�[��DTY������/fH�|�pr^J�,E��\�/�����N����n���۫mō��Ϳ�D�U�c�TRĿ�r��~j�FR�w%fH�c���m�A	�}�
����$����/b�y����F}c��aW=X�i�?��:�y�7����g�'i�M�wF��r�.'��}�y���o�sT�Gy;��;C+��ρj�2r�
�Z��C�	��N�hqJrRU�YŬd��I� �@��A�۝-jgIpv��R��S��Z���gB;�c��*�ϣtٕ��	+]Up�$P�b���Ʀ=�3Nh҉����g5���S�21%]X����<���D��i	a�c`�*j�>zI�.-���I��C�Rs�+K�|
����,�Nc���AF�b�.���X�~8��z�X���7�T�\�p�2%�}���'��H�.�9�H�^D4�X���"Ȣ��T8ڒ���Lm��b�~u���w&��r��r#�Q_i~��޷�j\���B��LY��>A�`���.�'�r#�+R*B�/�r�K}60�`��M�D�~������W�(	��}D�Jx�+L�&�n=�-��G[m�xs�xU��`.!�*0�9���1�@��/�S#f��D�$�S��oHR�Yf�n}Y��À�6�F� ��DV�a)��5b�J+�Q�w�0���NM|��.�����a�="��,�����{0^j?�d��[�Jўy�iAY�]���w�*�r��]UMc(������� NnOE�5�W�{Iiz ��lJ�]�$�ט�4^J��ҤX:��۬��L�ғp٤%r��mSg��y<eG ���e�"y���Mr��$ȅ?�3��K�,����8�+yķF`n�0�(�^,��!-��4�:�QxHz#�P����/=�V��ڍ6�.\K.�����A���S=�7���&oAo��4;<�,�}��8��W�j�x�}�7T�����պ�b�i0�#(z7�-S/#�7FC9X�PH#C)�/J֦�<vFp|(Ț>�r��׃��4J��A��Ȍ/�+�M��A�i�@*��R��
i���S?%`�qhs����\�k���bd��^F�!�N��ѸB
�L}V�G���s
��@�91h��D�=cOo!R&ExU��z8�4o,�n���e���^0�C� y�hp�^ZOݚ8�_m	�&����1��W����;
8$�p�JÁGC�=gp���,o�>��#�Z��F�&I�j_ER�`���MB���1R(|��.{����ls49�Q/}�e���IXm�<!�����]F6;�^&�}Y���v}��d�E~s�������u܏
p3���Ȳ.,��Lr�<*#J��644��ȳ���+y�B�%������:$EJ�!�b��*ad �t�/��Ǭ�.2��XD��c3֌�
���l��S�
�1<�v"�v����f�,���g�8Ֆ-���Ƨ���4jqA�? �ФQ�F�]4ws#Sp.�3t4�j�Suⶄ�8a�ONj����qޚ`0s�ڇ��=��f�f4�\����;�=����ؓ�f�m;z5�2�+S��t�֕�P}X3 P�Ȩ��ց\rDs���@�>��� It��!�p�?C��ʫޡ�"�d0� ���w1�Ĭp+���D2�w�q�;���"Yo+�u��=�I�
� KAi ��|D�+A�n)>J�Yf���:Y˻V�Лm7OX>�逢���'/�X�V�������&�����1�]C�z�JC�8�o��qI~��Sp��0����V�h$��W���1��vI&��f{0&ڨ0�rG71�r��RK�v<���M]#�)�a`����!��g[a�fm�/ּi��:lMe4m-1s��Yr ֪��X$����k�}v	��qM�����N����U�� �2�����T�\!���I a�T��g��B/���d���ϋdٞ��[���?=��8ػ��y@HPwį4��;J;V��T����*2����s�%����)�C�Xߚ�VrKod-&�z�C�&��n^F�G3K!�گ��VJ���og�O#z�D�uKt�'f�	ѴN�Js,�$���t*f��B[��U��_Ǻ��������`-���C�X��"'О�=�8���`������v��Y���$ϸZg�T_^�܄� ����\��ڲ�ʬ�>��Wo���}_}�����~Ro�lR�<�=]�e����_a����G������q���:��!�����;�Q��������b���O�E	�b�E4zr$�ׅ��]BW�P��
@�t�S@ƕ�^��XR�X�_K�)
�!���7���xI]_~Ei�%H�*#���b�zi+)�a��]�]&I������+�?�5s_Fu�_��0/ٝr�����o�-��h�҆C1��س�:F^�z�V��������RuS��+c>w�IN�dN'񁜴ve>� V�{!]8�O0A�ԛ.�;c���WgI�%\1P�Y�f�5�N�|/�6k0¡4E[�bޫ�oxӔ*d�=OG�O���;:��#���D�~UCO���	�_���"YZ� �8��y�A�������|A2�j��WQ��˞G�6ͶhfU�$$�`eC<�U�,����$�n��|������i:^4Y�Y�Y�l`b$�'��O��Vb�L��R�#İ�2v�Gj��*L�#����ɻX�&�J%E����MA+d��Vj��v�b��GYj(��1�I��C�u}k/�a�f$�Fᐆwm�I0hԻ͋&�t7�k-D�y|�xUM���ވ�ױ#�"��e�4/��|��Q��C����v�K��D�Sӱk�qK�Ck�k
���n��[�����%)��`H���(#�=S|O2}[ÖK�f����<4zC$\ ��@�fp�&L�a���5�:��ɵ���tU|�ޭ��l45qߜ$QU�X�[��3�f�3��®G`��[��8��D1
4�q����-ުW{+,��uU��|=�����f��G?pĊ�)�C?K������8���!h���1��H7th��u�j`RH<I|p=R2g|�g���;5c��ĦK ��x�W��L(�ċ��� Q"�Y`�ʤ_"<���>�P��~�E�K�WX`��8Ašes�s��f��{�t%��^����<:b�k|�U�(�
�{ıq��VW(����Vj�J�O���u4��2����-�${ș�K{�5��)��N�c����p�����v��)�7"�ݱ���	I�:����t����ފ�0����+�����G]���\��B4Yߖ�?��&T� =��Ŏ��W�J���1�����O�j���ɛ��(Q�F�0�wx��|8�?�m1'ӛ�3�`/����P!(1ݜkB#=5�*2(��k'{ 7�̋^Y�TП�sy��B鐅]H�g�\pDCM���2GF��#����ذ��*]=����S��x����ב`�f���g"=3̋�
�>�����C���\G� Ye���K��@��h�LG̏�0i|V��_>�U�m���=�Ϡ��tz�*9���ʽ�xs��HEMo����>��0Jj�"GX�\Q�Ǐ݀������MZs�¥WĄ��+o�����R���Ab �@D�-���k�JQ�?�LP�Ո.�z��[/�D˳K��@ڼ�:N�.�u�w����a��ɿ��D�{R��ca��lvw�a=��&�"��i
�r5Dŏ�r�
�ƙ��	٠�>a�k�Kxcpa�o}z��>�=Ӆ�ƶ���b�
X�8�n���ݦO�Wf��$Vo�,3Z*#^��rh��K=�붾\�F��V�Xt�6|�����0s1DO�xOߗ�Kˎ&� �J%��ź�p1.उD7bUf\��=H�쵹�nј��]������"�ͺ,������b�����aY�V�.n�Cin7���"���vj_%D��A��ՐO�`�c�yQ�����{W8v�{�B���u�ܵp���sM䙺��I�Pi�B��mi�6�BW�X��W���B}O"��D�"޷�t��a�fy�;qp���jCAg7��O�t��[$���XOq�8��h�->���&6�����D�͈���~����U�M��{Ua~r5$t�21r��=�����:|c��:<�g�u�y>Lm���\w"�aZ�Ybсk���*Q��202��e�HK�!�be�HR�� ���@��*\9M���؞M��L�����W��<[�ٻêIA(ݓh�Mڊ��I��C��Ūu�E	p��H>�s��Ͷ�[9Q@F������o�bíH��$��/�����]"/3z��������\r%�Yt�Ͳ��|dx;�\E����o���2�����У��\�(A����h����U�FH��{kT�_ˏ��>��\��3���лU�Ǆ�w+8���� ��"�#R��6�����)0~������R��s|p�"�r��v�׈��Ύ��o��;7e��3�_�qqr�]������{4%�I�Y芗į6��bHr��㞝i�o�N����҆^��<���"荡��5�j!x��<D��ޑ��[�T��C,8���9;Ah���d����=OhV#�ꃦ6.�$�p��rbT�,��(\q/ZC)a���xv��}�kN[T�m���~�J����o(i��yc;?k�˓�ԃ�[o�UvDЏn�b�B��p:�2����"�+u5�nS����W�%��Ie�ŻV��R"/v�i��!�4>��#�I}��&|gjO�㪆B-l^Q3Pu	G�-�rg�=����K����I0�YE���K�����5�)��7g��xQ�p4)g��5O��\��Jv8*>Ϩ���'�1�	�r�ىbՖkX��,=�I�ROv��0��E�r�u�g���|9����TN)q.�l�����!���=0<ֹ*@�e��P�����c~��IKK/�S<�z{���]�϶"��d�J�!����%+���z6�I�U�Jr�F��2%�K���B"l�~
�ҕ�4)�6�>	���pX���Y��q�A�k���@�/��#[Nz6:q�i6���Ѹ�6);t��z�q�p��c��������m�-�k��J���z����'�A�&���]ʠ0��N��F�=?���lP��B��-��o,��T8<���7!��rim@İ<�����e���+sHx}(f�9��M���[�[�?b���=����g"��.�Lji�E#���x����.��oR�Nl1&����Z��	���p䙭>ͺ��Ǵ]$���M�q�Y׆*��aT)d++���.�������9�8d�������4 Ҳ9Ê3�iF��♡��@���6�a��S=)v�́��p�m���I���=�@;3���������*�Go���4�@͠����:t^��\Mq�x��a�m�5T�t��-��գ�S��� ��GH?���}�g��*�(R��(IA�� r<z�hD�F+	m)���.�rF?��M���HM��� F����7�+Q��Wk��I�Y���sա�}�Q֪.�$"Ƕ�[w�o�qv�YQ>Q������W�0���Z���>rں�x~�Z?��ձ��TA�H���A�4��.їH\�m��K�|��9X����C~^�#�X؋,��˒$S�o�������n��V����c�4�.���X��>L���F}m�Ց�n�Ϡ(�K�Mp\쿘�1/�����J�[�����Ai�)�#���]�@ٹ��:�Ѓ7��>�(��%�S�KC5DZ蒟⒇>1���J$��~���e䳂a��y"������ϔ��uXU6ļ�B*	x"̱Z�2�-ܸ5��s�5�q�M�Kyh=�iަ�x���}m�(jחMp���n��Q\6^�/�a�����K$����^�X�v5M����S�?��OX�8�8'�,4��,=v��+�o�-I�O��������1�*��+A!P�%���ǀBm�('R��p�H�aX/N�H��b)�d
�q��~�Q�[�(:;���׆���d%�n�1<	�*���ǵ��C�2c�����sd��ԅ�}N��#i��+�qt��?�s����M
�3�X.�{��Knz_(��@�K��+�yޮD��7�HI�C�gy��{�UNI�MS�Z���Ӻ�����Z�����1�h���h�1jN|%-Mċ7?M�|U��Rs�f�'��� !���{��A����5W����s��U/� )�c�cX{i:Xp�Ґ����)�j� ��q�̈�u�	e�A�Y%��ۨN��J!¢�t�h��D�` /IB#��� �z�|��CD�M	G�[���ˁfV�6s��� �7)�%Z����x"��(��l����h��(�olޑi�I<��.��~���Jή�Y�߹v��x#�l��ui��̣SE�@��q����2+�4�i������jڠ6cT]h���0&���骤L�{!��! 2�]z3�-����:.fgt���"|��͔��L%�O�(ynl
�u��g��|͎�͝'9�_�yDD�eVtV�>�aeL�O��a�p�.,�sY]�������׶��B���C0
UR4�	�Έ��C����:@�g��Ӥ�$�����QpDW�t���(y����^D��8���{�g��35j�h��3�#I�������&�u�@\����ݭ�,�,�� d�\-���]��z\r�f|�K��H�>r�f3n���k[�S���>1 ]��w�NU�K��ܔ8����C�|����\�->-���O�Tb U��A��1�pP�;y!� 
�p����0#<���m�����!g�Rך�Zh԰��1�<�	��yk=_8HAث>kB���}b iRP��ߞ���L�p�44~*��Q�
`�Nu��1c��Ti�ڵ����Ȣt�9�O
�/��5|��l�#CY��,4�dV^�$V��C'��C���rw�<��i���n�#�O��֩}�J�^'�e���)J44��>-A��!b�4��*[�?]W���-L"+��y��F[+����*�5������C~]�$���7����:Wʎ��Za'�s0���:L[��Tm���q&Uh��fϞ�&�o���n�RvE�%�0ƴ�%1��o�!���k����ʍf����k"�,̏��#ݜ$�8K����Y�n��+�4�r�I�����m����r��R^�Pڅ"�ygݨ�VvH}�8r��Ԟ=e?���o��'�-`t��2�&���=�H]���k<��/B����u�@OpsS��'���?����?�:�Üh'�Gn�~#BYh�/ 3��)I+D'�����6��8!�I �'ܻ>�S����'h�m��l��`F�����oBQ\��I�	���&��О����"�����6��V<\ ��đ��N��;V�������8���A��ķ&I1�[e��}�;���SA��RoU��O�e���2 �L!̴�Q��X��U��MAp�#�R[-�􋻙'l����o�n]�}��x<]���ql�V@߇IP4��Z��.
�M�'_�e�-��67l
�M�fB"X]���i7��M�cB�|��d3�܇^��C*�NV@m��A]��:���W#��� c��ݙ��`g� `��s�@�u�T�k�Ӻi��@$>��<]�j�V��GF�MR_�F��yg��oiD	Zq�؛7�|�>�����BĄ���9�\��XT��A�+���`w��hj1�QS�P�FS�x�./SR��E��!)�:��
�ĖZbAeN�zs�]G!��R	ow$�������Bc��0)vψ�8�T��B���.���B�/7�N��3aV�Ӫ��g9Vף�I�[����˝�ġ���DO���?����U3�F��D����JX>I8�}�l7�����ʵ�EN0Z��M�
:Ss���d�"�0
ک�.ӨA��F\s���%"%�������O\+�+��b������*E8��(:�ȧn�hЍr�F}t��z�E�wR;��Ev^��������d����!�z��"2�tO]	 �����]�Z� ~���H����%q\�N�|6�Lٵ͞^���-�ϴ�he�����e��������Y��V@�ٮ�0)�4̅�H!�M{�2�EG 6�.͘�/�:�Y��:2��$�Ob2+��P ̿GUû�%��md�ʀ�1�ycCȪ/�F'�a��[Q:p����\4��D`I�{��b�D}9�n 6�� 9I��_���=��c�IZ~I�Y�m^�Za:f�����o	�Lu �~x�bp7�3�g r˭M]6f��%]n촲R�	�j��d��k���
����C����;��G�O㎋�����
#��k̯�ڒI��2���z���Fa����V��a�.)�o`�����@&,FA#�[:�O�i����f����$r��d�>�jU�7m��@(o����ua�ֽ��z��3�!FrK�4|�)�GK�^aA⮶�>�}T]d=���܉����wv�l���P`�-�\};��J��f�z�Q��qr�:G�h�ŏ�	��L`�nn��v��Z���S����W�!w\i_�����0��>����E���;��*�[�N�X�`N_�I�)Ȇ��3,^�eC�*6_eW�
���%��;��?S��܀�ڎ}f�;㈊���m��:�B�tp�9�k��� $�\fY�8%��Ǘ�xkjr���~G;��r�f����,:�t��KR��ӱZ�+����?�'�y��Mٗ�`�"�Ty~�����%��weՙ��`�g�23
Hm��(I�C�DT)�u	ţ�D�,��y!%+�Z�hL�T[�6���W<�	h��hżVx��>�<����a$�|.×�'Gt�@��ys��/ -ᗭJ��l�#�v�S���-�v�)���s�/k�=�7�~wT�9FhH�Ih_���tyX]����R��ͩ,�ShQE�qi�7�ly2���0�_󢠵'Z�!�.wZl5:u�l�E�+�w!l�Ƃm�#�����`6�G1��<�"�c��t�̍�ZćnIq�C��iEm��cR�X�R�-���:rrJ���\䆳c1`��/(wws\p8FDT_�0ˢ���2k��wD���Q:c��n���O��-l�W���G%����k/��m/����*�p��g��ƀn����p�K0"�S�q[W���6 ȥ���|�L��po��D��A!�x���4���|�)�U]!ۓ�J��	L�謺��7��O�A�xt�8S�x�G��l����K5ux����S�,$j�n�Not�K��ɽ3���f�x܋N
��h@?�B/�2��މ�l��5	�if�Fn�F�����	�bޯt1�\ig�k�K ����uډ��3l��Q�H�r�<��d9�fJbU$�T��˖��1z̴�E�.ډ
�D6�<�w�M�����K�d/��T��z"N�xSF}:ض6�v�ԕ�+���`���M��N�q�_��%p��O��竾FiеB�Bl��8���ȓq��H~-~cz6}v椊�B$��)����,Q����L��UEzwy�����7�/sJ-�SE?H���`k���#C�%]
bE	��VA�Q�Tz��A�L��!6喹�lo��l^������l�bro�9P�q�`�cx�y��z�I�����#"��kb�-�k�+� ����՞���:m��lǹd��g���ķ��M��ltˮQٓ�iD;icDRJQ��ڎ�3in����`>U���iL�yw��+��\�jgJ���{�%B;�}����/��=j��m<���.��P�r��
�XcV�(el�$GZ�_'+p�NR-��/$�9��#-��V�6l�֯M\���Go8{5��� ���������x~%�Z����9	Ʀ��v^}>s|MG�H��7������+ϼ=�>��	%f���je#�y���5{�N�[��Č��;�J���(-~�S��5v�G���2]�EHTS]?D���He$@ڊ}wP@���t����l�g��ݤ���-�u�z/˰8�W���K"$f[i�Բ0De7ѥ\��ݾM�;���PW����E��5P�i�����q�+������bY�r��S�*�J��˟CC��sYh�6��oխ/D˾[���Oӈos	Nf�V�٣�����A��#5�k�X(�1�eQ��[o~�8?Ӡˈ�s��1�R,�W���
SI&��{�\tP��
%S5���)���b���"�G
s��W\>ۊ|��S��X;�˃��Om������p�wQ���_�;Ȳq���������8��Jux+x�@q{�h�'�2�& M�)Ǉ#�ɹ�c��������n�
���έY�)�����Ƣ,�VQ�j��&YMvh��]�����!\@!}Yj���;yx��`̻�J�zT���u�z����wD`��mmߺ2ǏR@'^԰���o�Ġ'�o�c3���i�}gw�ჟ18d�.Ib�T�	/�_R�")������K��̱��3����܀�t�:����V���_Un�y�߀ޭ����.Y�3p��gB�Y����E���7�Q�!t�AUZ�`�e�j�xʑ�.�5�{�Qٞ2��m)�������҉�5d��@K]RO�EG��z&�[}^Mh��)hm�<u�!n9�ņ�a�5)�kL�*���� �Fj$���W���˓��<i���d0NՏ�<3h�Y���Xb�����+�0R!	����I����zz!��E�Z��/��5��ps�a3��)��C�,տ�h�co��#`S�P�$�.����EX�7y�|}&�U��O�_�i��^b)�\-�[�O.�"�<q��U��Ʌ�h͚Z��u����pR?�A�x𩧶BD_�c�I5(�*��n^cg�L)� Ih�@�W��1�]� �ˀ���4?���Z�E�f�Ub���.4i��Б:M���<�,D&R�[BB�יqu�rɴ~��X��s�z�����>���jME�z>��_�Ý�J�8���K��el�_��Â���%>��r��:"�-ƘĽ�����I�������\|v�қQ]/�����.+F��n����R��H���ׂ�[�G�5v
�i��*�f�}����7��{ �+�h��i��̇ &�JF©G�؇)|�[7V��%��$r���d�A�O��f��N�=&Ԝ�v?�m	@Z�=(\�����c�i~��of���,�7��*�'�4�"Ff1�+�+�["<���ߐ��b��W������,����=->�&as�Q�M+7��	��ɟ�{�<�FM���3�i��Ŀkm",@v<�`���*���l��{�	��B<�I)�M��]77� ��h f�M��������HQ�"gY�N"�V˶s��۳2{������E���VIl57�"��Ր�ܹH�W	MB����;���Y�"�bǶ^�
�����o4����{�wo�� f>I� .���ft���H��Y�:��D�\��Ԅ}�hB[�s�_X�ɼS���=4�?lƀ�v�|28����4L��=� ����S�z�6��i����5�Q��Z��-�8h����_�h�h�Rć��39�A�W��u�5�*�<(��-n����=�k,�z�+���n�����$	����(�K������y��1�'-E|��\�X(��:��*���&~����7�OT��m�l$�c��\��3ē*�L%��H�s���:������Mh.H���Ұ~s��-=�y��'6_��څi��T$�v��ݠ� ֮9���p���Q4os�;$�%��|~o%��\�O�{����T��GA�V� ����Q�r��`�ᇬ'��c)�D��@�Lh'�`�ט�`T���YK����5�+JB�q�򔺓XK�d�M�ܸ@�*2���_sc\��+��@�p�<P���Ҁ�n�KNҚ<������eq�����
�.0["�V�)��״ô\9Ԩ���^��xߖρv���R��c��VY��_��.��j��/�A��4a-e�MPo�n	�+xM����g�4�+��)Ctd'�L����a2a([bc�FX����kՁN��2��M���iR����`r�c;c��<~nLˎ�iӼnKE���������*\"����C-P<N���|o2(�W��{"lA	�k�=G÷u}���Pӧ�*���E(�_Y�s�-��h����Vt-ZV7�+"�\ j+����U�0�W�+�'F�:�X	�4��2�V
D��I4��/	� �zn3����O|u��_��b5DdH�_|</�`-؄�}8,�T{���g�+ƛ���G��0I!C�j���j��c_d]J)�b�q5q��J菗+�o���K��� �泲r��^�m��~���66���Q,C�����΂	�W����?��lFpVDQ�JMg%�c�AF7s�y[�]�og��n�V�aɪ*�� �@��n���^���5z`�Gy�6��>x?���Æ�#$b����= Йs��	S��� �������4G�'�	����vJ]ˎ����2(�.�����[.y�j%y��~�ޣOկ|���g�Ѹ���y�FdD���/2.�ަ�j�)�%��r��.��J}Á�H�����k��c�\/��ۃ�
|NӤ߮�,gM�B)��Lv�M�;�B)��Y��?�}KA�j>,Z[m	�	�YPe	2(��.H�4ť��6|���Ͽ��T���=�Q�;f|��hCz\:ū�������J3v+0D��_#
�Ŋڀi� ����}�g,��dL-&�":�i��v�6�r���ak�	����1����\�~�2��ag:{��w�K�j�V#��X�]t�����ZJK5Z[1`G�@���B<���5aA�EY�'`V�s*�4��C�=��
�y ]䧣0fP���֭��c���f5D{f(I0�lU"����&/�����g����CJ���R����u�C6u���15:��N�}�e����o&�֥C.��)X�B��"7BXd}�*��k���8����bLyKc�l��[�<�OT_�D&e�M�N0��"ߤ7��jQd��Պ���l�d�XO��Q�g��bk�ox_���Ҹ�0`�F� ��o�
�E�k����x:��K�6=e��J�����_��C���hz������ݢj��S���>�����g7"@ �S�t(_D�ep,Ԫn.��7�a�Ⱦ4��V�+B�]jd�?�j5��/�3��L�v��md�器U�OR>�N�tEhc(�S�����<�mv�&i`��D�/`����K��vBz20l����B��_�(a�'1<�%@9����ć��/j�$)*<Ǫa��O���g-�3��ǊR�q[i���Al�7�[��>ɩB��T�j�h�K9�\F���=h@���~g�
����4?k�e�A���dp�̵ �=Y3pg��_݌ZD"h_/���ñ��i���&�>��д ��M�RT��_{�ѓ�L"�+�,�?���� F��2GB�~�#@*K|�;F|(�Y���=c��: T�/�4���zu~��ۮ^��埋�~�ed�B���ؤ��3�6xK>ʫ~�:����ңJ�r4򆗥 �F��8�}q�Om�ܨ�@%��� ����)<Oe�3��Zp��p%%�z^�f�b�0 �U��uF�\�ċƉ\=�en��:�.��W���ڎ���M�Ԙ�Ch��H��7�	U�B5�
�������fr6���l\�9q�t*��`��K|����f�޺�RB�������#!�*"5�
�R󟓅О�6@�u��N7�R�0��'��P��؏��� 8�����|?�@3��Q�&��M�52=�b��Ţy	:��\���
�dyY�`G30Fv�6Gy�C-�{9�V���k�n<o2S��Kw4ľ�zc�Q�{5G'|5WCS�g�a��^kF��޻U�b����+�x�Ɂ@3���1lS"�]c-����לu��n���x��D����~��9�d���dxl��d�Ef�X��W8�;��o���=�L�f&��62�<�-����;ʁ��L�W�GOp@�C�U$d�r�% )�@�1-X�
55�Ǫ�04<��0��kz}�m7���Լ��PJ�t%ɜ3e1 �6=y�^�5 �X���L}f� �"(��c��A��5�� d���7�������r��;�u�"��-�qH�.*����o��놝Z�9��M(Q�Y��Ygb��B�Q��E?k�Os��Ŧ	��?��e�<�@(^/|3��a1^e��1B+7R��w�];�*������nE���9�gd�G��,�nm�KyL&���b����`�7���ѓ�ӜkZ�V���_�O�����	��w��z�	R�r�a� O[���Z�=�;�W�!7&�1��E�]:"��]�\���E"2C*n5<�8/^�5�v��jD���F�v�������Z�&�r�lj2�n����I>��W
�cρe"/g̹��7_���<�C��\��_ȶ�<�L�O�ܪ�D��G.y1����w������sZ/ͤSf���<��E���?g�YG�Ri�h�牆�q� �@,Ϟ@����wI:������������-�K���^�ս{1Z��>�v�q̻e�5��<�b����SO��O4��Hؐ,�K��ӎ;Zc ���_�%��G�7�!�&�}��7N��~����5c'~~���Fǻ��=s��V��#�,��w�� 4�I?v�;g��&��}h5E��wmv����)`T�H�er{���Ϣ�y�U#�������en2��"���1٨E�_�V����{`��M�j��]/��Os�^�C��r�i�@>%w7�ވ�BIcOEs�d'-�����OBԅ�qRu�[����_bf7iW+5���YO���D�����!��l<��d�q�� ��z������K8J����|��_�����o�၀.26�B�S�����J^�7�+��~J������Xe�$/y>���G�<.�l�::^��c�-m)&����������"s���P+I. ����ՠ؛�"%0��$B1�,n�VP�.J��2;-ᄃ���28s���%�T�m�e��b�+���!n;��zV�`Iu�0hƕ��K�r��;���h����'�	vdI�����D�m։)�� �l)0�����#�c鼶li{~�׎�X�����.N�P�$���r)�ܨ�ޖ|P� ���$i��IӁq�r��~�&�e{-\:C��D��\�Y
�R�h��+�2<��P��+@Mq��tW������+e��h�#�վp9��pݣH"��eJQ������ɺ��cJ����|�ߕ74�h�~&�@kD�ݎitBi*Gq�\��Vp)���J��+C����yn���f���e@<��S6�H�>(��'#=P
�i���zc��B(�t����iMi��i�@R�G��lO�dT���q�����?^9s
K��cl�i'm��M^��Ru1��Yn��-Ϲ���d�>���y$���h��ٕ�V\�i��%�E
�c@Dk,�W�Vc�t8�D���d�Тޥ^��-悈3��"h�)^j\I�Kk�
��R��)�Vš��=x���hBR �R�^x!h9Y�B;��m��c���e*.\��Gߋ�W1Ú���[#sц���LO{0��n�A��vHe���u61g,�s�X�ux/�����𿛧Z��L��N���vb�T���� `�}Ξ�t0sMo%�Ar���:s��&y�A[Z���r�׍^��,�/�u�/:�G:�@BX��X��`�����V߆h�νbE����b9M�`�ug���X�^W���l��-�����^���)��P=Z�0��R��Q/����C���h����wG��3���D��i�Hi�TxG{��I���:��^
�TV�X K}nw8����R@R��jj�.s�׎���˲�"ҫ3E�o��͐A�ЛOD�%���qH*�/��]y����j#Ȥ�EX�Gi� �e�ݽ%�O�����R&r�V/8�7�Բ������)E ]dG��T�.�uXT֬&6�͝ypiQB��Ҽ�\����D@/�~���p�Q �v�*Z����o�c-��6����h�GI���m�GM�N�a7�iG�J|\	�'p�U����a��g�e��)�t��̢�F��cwN��ju��Վ�NV��BN�E�g���R�.Zk��BM��x�ց��}q3&`���vP��x��$��w2�fեf�����N�^C�Ǐi��E���G{���_z2׬����!�ao=�8�q����I��w���8��������7���;b��A{o�������Q��Vs/���)�K����m��v
-�&U��?��b�eC��a.>����v�ih!eܻ��h��P檞�(�Z:��}����JT��� tzj�D�*G3H��J�u��`���xȞޗ\oS�o�8�>�d��4Ћ�n��w����J#����,��|}��#�"��zY�0;���r�-TZ�lb͇��M�4�Y�=T��i=�؋ӝ���|�s�ՑV��D�1��f��n6{Ϫt��vD�����@�A,z����q˕V���i���g/�pO�1�Xf"4������gA����>�g�^#����%&���b�ʨ�NQKu+��G� ����LjS��	��>�� ���Kd��m���;�������d���<w��c�����J�NNH>Ę��JyU`�I��V��ѡ ����Í>R\�s�bCo����ѕ�<���&]q�;�
\�|��ϭ�9^�a.�6
�/��"m��E�Qb�=q�٣n�M+�R��ҍn�&���Yx)�Q����ZR�u��{��@�- �:(|�ӫ{O��������>���ټ�a��#$`���7�I�������E��?��%�[>,���4����+~MU� �]��R?��]T$m���̬�ʀ;����E�,}!������ѣU����el��a��_�=�����*�,��� Υ�7tQS'.�F�}���4�O0�~�1��քk�aw���X��Q��9h,��uF��W�c�P�����p��	�h���C*���F��Q�'ٱGo���n����tr l���iW��:��"QƘ	��D��o�0ä�/6I�0o?E�k v2Ϲ�+�\Y��2�"ۖ�h���mM�Dj�*��3��"l��W��AU��K��:V4:����x`�sHsUYf�)"��,\��		������,��d�� $�x9<�.J\f���^[�dUv��tc؀r���?�+(V�"�H���'��f���/�d4��	�<��B�2B�j[xL�?�n�x� �vi�JΘ�7�q���|%2��H�5���0��@�e�'egO���57K5�S�հ<�ܔ���E��.(t
�u�a|�u0I�\\�6XI�k䮺�I��L)��M��X�Ș�B �R���#
0�P�����ʂ��6�~P� 9W@�\^�߿�li6 �&�ԫ熟v��!�;��LY�P��?�X�m����� I�:_s����� {���ٯi�Vy�~']������r�x���5���j��D*��ɻ��f��L�}�[�]W%���h$������i�>A·t!
��9�pF���� �1�o�������'����k��3>$R��o%W�D���["xF /gn1p����qU�Y��U��B�)�����n8���D��#�)���뗉��o���n��q�ɵYl�<H��q���AO�6���v��h�2�J�u�:[*+��9��-s�[*'�a�'��= i~0@�!�ԑ���-f�(�[��d��� ق��b+Q�{ZM��%��{ ���� |Q=>��>j<X�Ɉ[`�)�tz��e�\8�?�#���38�5�
���� aݻg7Zn�9;=^�F��ߠZ.�fC<r�t����9��J T|���i��̎�vk��|K����&��`��e)f�hUi�><����L(W��[r[�Y
�p�AiA
�"��<B$}�ٛO��֛w0�O6_�ҽz��6D�DTr����^��@��;�7&!^@� xټ#2��|�s���6�����J�GPa�7����^�lZ�k�c�Y����ΣiS)v���d�N0�u�$��ab_X;�ݜ/�w��oA�'r�B� xh+�2��ij?OM�%�sc�4�7g�a��"_��D\�����j���4�1�U��j�IP
�g��N �0i�"���ɒ#�1Y�R�HDv�|�R��d����/��Y��Y�&���-`c�0x��p0��3�M<n�#L�{��3�d����H�7�u<S�GP%~�}�ƨ����e��5�����3�}3v!1����e1�S�:���'ޫ��南�dir:��=M�(jO���\o�������E�)�n$�͢�Zp��V4
�XLo9
�v��H��{�/Z�d��C���?�2ѧ<���W\}Y�TO�K	�3H�Ze� S6����k�Uם܇6[74 �pʢ{Z��&1e��bV�����_�T}�-s'O�P>�u/��.�S=�$�Gz�r$�����R����8'l��͟-�����o>-�3%|0�d�~�W�*��nv�bk�=�Dȯ�2`J8��Zg2��yӸF=,��j�7�?e���N�H\��c�6K0�^�Z0����:S�2��|�F TS��\3����{b��:�Ka�/�P��ݗa%+t�8��1+���Y%��*3A����퍒�({��I�b��Qr��on��/���+_���ĬиT�]���e��R'�1)M�b/@9��Ct8�&�1�K&b��q���x��1qNR��m^�1�U�W0������[��-�:iv� *Y1�uSod�z	�[����!�a:��c7�E�UDZf2���BCa���QW�hb{����_Iݹ}���Ҩ�.�˂ސ�"��I��I@f��lYE�HSNZM��'vS<���)V�^M�yƐj_<�ֽ��#�s|���ӂ�r��6���0|��"�1�4{s=)|5�g�����!�@n����3�u�~�kZ��T�5oDg�I�F���S������9���A�����u*j���|��l'��Iy�*.�4�@I=����Q���<�Ay����d��}�b�4>_���$�߾@	�������13isί^��_�;]t&��^��ޜ�o��lS�B��(��o����EI�)+��0��FF K��P��8um9%Y����şpC[���oҝIu�m�����5G���A���1�	z����8�R��d��j�a�F�����)ɸ(E?,��r�,�Ƞs����1��*^��;���$$�����Y�ב�!8�%���N�����_ �����𻗴�xV|�)Z��k�wj�)D�u#WD�U�I���@�ƞ�¢0A���6���Z��>J�)�F|�k��j�B���Zh�$\�C���7SR���7�F��-�Ԙ�4����0j�x�ޱ�n��W/�¥�����+�zF�5��M�Pzt�;7ī@a�o1s�	k���1�B��X|@�&�/b�pQ�Khւێ�L�3�Xs��%�� �X����Î��S��R����_b�ױ�����6t���H� D	�M�YoX������6{���%��̑���\?B&<�K� ����H����b�5����秬�7������G���K#x�f'�8��=��I[���{,q0�M�	j��b�W��P�c[�PZ)}����<~�����q��7�{��,�D�e�*�H!U\�>�[�⎐1�@�b6�Hi�~�0���� ��`�2.Ĺ��PF�n��ܑ��G ��Ta�`;d�B�SR?��ǫ㆜�b�ԍ�%������(w��B
'��}d錡�����*�٠��T����@������
ٍ�]C�����E#��%Դ�͕�w�R��D�{$jQ�O����ڽt^���2\��N��� �����.u����������4�n�`U�5%����࿹1a���@�H����b\���v�gi�����Zٯ��C#URK�=9���|���e�| `�{pfe���f�b��O��
ܰ���u��؝�Q]?m����$ȅ|�!�^�@o��GJ���"$�b���H��"���z-�Ɠ-F�!s�-�ԡ�qRW��58�pP�uUxA4?���z��S����(���&��e�Lڭ�J;���Fh4���p=��C��R<`ky�K7��
��4�����pa�>8�W�ކ��y}�ޠ,�3û$��:c�~o�����N(ev��nO��-�d��G�N�e8d��~eR�ܧUg���=�o��)t�P ��w¤��2�'��s�O�L=Ϋ�^ӑ�k�;*pA�6yʅ���w#?綵t:ws��-�f�j�h�p�n��KS9�zFЂC%�R>�}F�E�X���ʭP���	��� �i#�X��%�Ζ���Iz��Ǎ�fP����l ��3ǻl?�ӑ~��'����"zoĐ'֛�{n��H�!47ap �/�㎫փ=9��頛��Em1dq��.aw ՔٕT��e<�F�o��'��>�גz��tY�<�A-��ϲ^��d�����w�x�r���2�rδ����Bɭ�y���M�ܢ�NI�������NKN=Ј%�_)���*�
���
T1���]#R˃��:����0���+q>Jf���`�>��w���:A>���*xk�m�6�����%���w���xy�j��9��I��u�s��MI ��}��6"P��%�����+�_~�q엱"�k�R�i����Y	�٥X]2�'Yg�21oC���ڀ�T��@�]�)m�<��+{́K!`����.����N�ZuA~B1���r�C����5ai��2�:��6g����.��p��#�L����Apb����������M�!neBuЛ}rPRr�4����q$|���[٥Z��S�6���e�$钁�ο+C��8rdf �p����KC����=�t��)��n�B���H���i������U���,e2�� $r��Zt�����&Mf#���v��s�s�,��iB�M�t�<u���G������$$��G�az�j_t��r���+�]�������$�P�7Yt���|xX=+KV&��)�+Zu����qIe����cn��s3;j�PL���`��P.a��?]9���Cs �4@S����rv�tCƙ���Ѫ����K0��#K�͗௣�ǡ(Wd}tO�N�W��Y�?�o7��&^'3�GG�E�mb@�IՔ���/?��K�f��α8�_"�Yj'&�A��iS�a�ʼ��
�Y$�8��q? �-wf�^N4�u��nLxԇ�H��m
%YV3��ʢ�7��	�+T5�1h~�r���:3�W2����/Kаi//��3$���.s�_�.�í��ͳ�Aw��Eu(�$%�X���H�޺W�%��\E#�rZg��(�I����!�����3""^4RA��Z�f�$A"��a��APeG�U��rP�WM���G���P��y�\�K���a;�gDلhJ��ɗh>���;�,�g�1��y�ƟÌ�;:)��o��4�9H' ��lL]T��@f���5���v4����`}�Յjq�ɣ.���x��&cw]�Nޔ���6���E�O_�2��ڡ�#g4$��c�a`��X�H��	�TXB�o,�U���*�vT�`�UᱬD��h������p�J�،�D�f�����yW\ut���V�&�!5�7^�[9`��*�J�\	����<f\|���5��*�5�g�s�=�!z�e��h��A%̀�!�jX�Oф}0{��be�JP��3��N��1+�O�-��T��O�8Q���������[��E��DYg��p
���܎�g���? �M$��]8�4�½�=R�,]�:��[�n��
*h�vo/<�+j�����h����;�^��g�P�TK�v^���$��B,��~��>}��U�p��j�h��۴�9}C*�(����Ď�ѓ�'���m)�&�A��p.K�y;�웶�8��S�X
3���=<�4�~�ࠔ=�B��Ʌ0�ꟳ�A�@������P[��f]��*.�㕍�fZ�]}RN��r>Ӯ���������7����E�*���)Kh��	FeG���,NwP�[<�81y��P�����2ץޞ��j4�+�y�k*6�)}�sr���#��<q���_�~��?�'4��N������v�a��g������?�6�������l��M���\
��*�5�q��%�,o��h_��6�6�@Zm[�r�BI�y�T���?vn�j,���� ����J��ućԃI��-��>9n��'��� ��6Ξ����]
�����G���F�,v�m ��f�$xn��9�Ë	$�z{��7��6q��b��<�ag羷�S-���_��X����KMB:�3�y.��;��V<8�D�/W0�sR�!��'�ޮqM$Q�Ԙ���U�
xy�Q�d!Z-��\��<�b��AtUn���]'��ʃ�a��~A��H��^�?�ם�lf��V�< ��|Be^_������ּ.��Z�F�G ��g�E�5+�����j���&~���G��3�Cؕf��ֻ:b�8#�
��MK5��[�C����}V|�*��j�VWo9�����[��/:�Ó����i�دOc���9lLG�����|�F�)+���={����t�ʎ[
I;��^4GS�G�.�{����J�mm�Ȍ�3ui(���e�kU"��e0ڭo�6��x�Hͽ�A��&&s��x�N�wܐ�d���q�-�D;�t`(�62ڂ
�`���1]?��d���(JTǜ>���+�Ϻ0��
����N���/�����'�a	�%�1�_w���&��C׿�+ ��GM�z�=w��iv�aQ��0��=�Q�$�?�>��q��L�e��2����$����֠R���`�WE}�죨iW�ͮ����`=g�@��.u!�8�+�6�$�rAt-e�����ѻ�>(��2�c����7!{�_��1�jA��{�3���[�l�_�;(}q�e�7�6lCgC�_�Q�߁�?|�B@G�+����77��*+������]�xA�Co���ĳ3��$x%�ق��n�ޙ�Zu|�����'֥�!T�X���]�S�l�;��R���>�Dm�bЃp=_�@	z)��<'�lv���*�1�yN�8EB�zD�c�}N��E��0��U�j��]��'�īa}�M퇌`����Czbo>1�8a�ˌί�<�h�9�L�zz�IV��H�}�����o�#2�45֊�zPȜ}*���? x6Rj\�䩶hf�DK��e���	1-�FewΘ����8;�ܮj��Mk|L�U�p�N9���49��xp��bz'�ݿ����M�Q�}�Zq�َ�Y�Q�"�(͠�HT�MN�O�������i�a'jsHd&�"~��>GY�����;ǒ{ms�e�ag{�%2�R�]OL�4g\ߚN�4���iא$�L�����	S�ܥu�T�0�u�^��#�ygm9,�͈n ?z�qʅ.�.|�X
|S8�
��oG��6�C�V���w#M!��G��̍��2  x��\�L>5z~�q���ɕ=�����вm��7o��̯��dk�r4�vJ���x�s
��a@9��X+<�8�ߑ�pu��9�H�̘S���1�3>	��-�+�b��� �9�*��X{��+��Sw�C�V�����Ԡ���srS�TQL
}2�g��צ�q�ќ��u}a>�-��q�*������~�@��%鱞�"���]�L����f�{��.�At/�^!5<H����2���O�4�Z����ؐ?��lj\�� �G�F"��׊&�
0���l�:5�29>S<>�|?��n�"��,�o�>�O[('Mm�2*��Rg�1�UY��}}�9�/ ���{��%?�m}]�9��'�#�Br��u�	�Ϫ�o�L���!U��5�S�Y�;5�v��g�`�L���D	��Hl���������A=�3���Ò�L�.t����s�!�q����/^1�sT�t�|G�y��KT�y�1���H��ߨ�g��2p2��Z� �D�����s1	���I�y�Q/C�Q;�N�2/�Ύ�Z�k"�7����_B��T�t96�I��a�>{���<&$��_v��m����r��TO��w���^'Â���Z��@���Z*Jo	Ծ����<�D�Q~Y��(Ʈ� �zl��EI[q�~���%��N'��6��11��w�H
��d<�ŀDT;�j�7 �ژ�#��q
��V��t�.<�7ί�	~�X\�R�a�_]�%F�1NY,@�D���$!.u�P�=2}�_-d�|0�����b��$�\���~��V��c�:ɻC�U���s����s��J�v��rmEj�/��Kʣ������lأ�F
f�x;k�����6�����F�_1�ɟ�-�m�|"�y����rAsl>+�: 	
FW��_�"�2�S8&��̷Af�C��h�[(]�q���ꅚ�Zb�'L�4	� ���'�N��r���j�L09��why�)$,��^mϺ���x�1�c��}�З�+O�Z�b��H��I���S�O��2`�I�K�n����=�{�S	Lڣ�ҋe�� #c��0Y�`�J�Q��b�<�@՘@�bzR�����激�3zF�̹���hi�o���+�/E���tN���$���fd8�;`	X�g��Z}���aa�!g�?���s�k��m�i38���_��A-?F/�-x�%��8Y�'=�$�U-��0��m	�a��n��-�J�AΒ?v��&_�+ජ�։�X+!l��k �Kkk*�R�J�����B�� �\��|�L[���T�#�~��-��؅u/�KJ�6&��t��}�BM*�W�JCl=�p����|yo�*��{���R��h�'�(�*�:{�b�<�2��=��Ķ�r_��F���T�Tuj�?�;)�����.1�,�
�����	f=��R[	�;��#�=�/�T�/�H�k�N窨N���E?AN"��g���k �{������d(S�Y���x��C��|�`9���e!!���,��!&*`��S�ӑ
s� '