// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Zh6eI6GoFL5c1Adge8vzeTCD1TtZk1KIzu0l6pBTqWaPDR3lBwxZvjvc7XtDzEZi2dCL3Dyfulya
PBtpY+Tfx7Ndjf4WjxWAwfzCOqY8sIuCEumQ1rhkNdiJBRBY2piQa5Fh+T7Ic9ExxCwHGARUodR3
MJ0w5x34vUzIMvb2E2EWIiXECEObOC8bH3JG8qlcSUjsQSRdgf0BvBTY88zhtcxEOmJEFsaE4+aN
DJveuccuA85GaLSzuuHjUuyHrKzaKWJTbLoT4CnpNVd0NN7EXsjHZHaZOu+1EhfJ8D65lxr+pcDW
uCniP4h1GdsPNzknbFslMMwQOnstgDBlAq0sPw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
0Ng71twGTtQnj4Y5Goe5pJPxKnNmS7Cm537GXIDUNTSvEiQqmty1UmXwej+JepMm0ueS3TmbjQxc
kFALUFrGNNLKO/cpJaOp6orxTcr93ubLRS7rNzGb6RaZ7/9UozxvvpaRyoPKwq98wSBqm3LErqaz
7q94VGzvurDG+O86W3OWD53zHYfg7ww35JT+WTvIKfnMU6Ka6kBju9jK8Sh0hZjzcLqHzBhqElGF
8SUtQVnuAAawo0QZyOBGTPPZOLQBxNeIewElhPYh/oe+khMA2Pyv8xs4A645vzbL0yOMxE5VeN19
NSS0sJ7vrtlUXLd1PbhYliEu9QIVEqNCgfIvldIVEGW4fNHe9Y/x/ED0rLl+rnwygUwtaufn1iNP
p0Tnim87Xa06DHoSl0EnomMdecOQeGOwtBuimOCdNVurVc+21x/jde6+jRwtENRVwtwYClMEREJa
ap+IuymMbxG5J0xLc4+8nwsVWx0iPsrSn0lhnA6sJB5qfca8tKaeCLhuDjYEfmVW+aiFekwwtDPm
hFC4Y2MiJVftLtD9ROuTSBp9SXdkzaVgV+TaIUxgfrFAwEQkzygkhAmuhj7k75MOEjgbsFBAGIAw
f/NeXFgNzuOMkf2nlO1JPimNEaEiREzN1fIXuUXxYAmstKrtSjf0JYRe2z435HScuwUuMKpFCkhb
lskGW6p3I7SOHzQ0dnHKbkKAlvJ/Xjn8Bu9S54bnSShJg33hkd5yL7yl1qLcYf2wkftqgiq7e9ES
cQbsEOohjJNfn2Q9npL+D7qjjpnqpIZ/Tj2ew6F/9DZqtpMTTX71pAKaLmKo/mWuiBULDe+dlgFs
nH2+IKP6iaw2ZY638f+t+uc6DIkG2hBLrQcVdmsy64TvIn9IanoBvhSfox37knFF4vREen1mMmZ/
XPr319efzP+d4SUcgBhMK/kQV1FmS+VddoL2of5rLsk+TuOSrQkZh6MGI302A6ymlxnixtyFSHvs
Ln2JxtwydlEMK4xR96D8RvaxzCeUj4vTXFAa7NiilSXR1A6tMhdl68MyQ5PgorLOzddEAty2bdZv
yHg78j2qk9lCGxMSKMqM2Izx6LSi2YkdvByu5MhKpWCPkHHJeqdSMVNZTjm89oJB6boZCH33cbWo
FOwJhCiwfOIXnjZof3LZyyoVWEPoDOhDj/ldD82c+1h3dge77LfT6yU6cp5LiXpyYXbVAWmaeFNj
m8wKfn3dCLrQ2oNFz3+S6IRqgWWqwsyxRt8bmKxXL3oVZnFh4NokBQv3tuFyaSrByQN3QZ3Sqkh9
5v+LaQdWJnQ/I5R022thNKQ1BY/welHtCzPl+0+H+Ed5ji+Tua5wD4hZhCO3Xd/0YS3y4tWu+ETc
yGm0UP75NA1EsvCgCQTp/0F9LI66Ffa2hE9EqeBEyVMWQC52kju6bFZjT7VWWHPMHKbYVNaQE+/J
/6gWrTKBv3Obhfp9sZKBMkctEzMJKlOB2WFtUXBaJCipJotSJVruRE6bTteOE/EPgX7K/KfSqn2s
K/ULaleMFEqLvv8OwMMJT1rQJ8o9ILmwQ1fFotyfVEVLuvDBni4FbnNBncnCee6qkXeJ35tZ/tTf
P1CLJOWFP9KCKfdds1ki9RoJs5dyk3eJpnVA/r8jwa6R8AhRUzc04pKRzZNcM7LbsHiG3TY4cER9
8euTDXich8GDlTbJxdAZfll3XI+StLjh3VGcBxa9HKhigFGV5OuZjjgnhbF+3GCawlsfsJsJ0ZAi
ohv/urUJReRu/34i83jWRcmd/mf4yVaVYnUSVxlaSL3IwYXdFE+WbRnDbph2+yE1RTKlnGAN2Oby
2xkq88XJc7kHDA8ueBlUiJmXoXsYUkDGRS5FLdbWtM32uUC7/B2HrpgVmgwFrSe5Kpoli6PHvdgm
MwfJkfozB2MlVa4Gx757VztawgeK1aagwDTeVZKYn0YbUsXtQk00Ciy0rfY+k8eDP62zAL46Ips3
3FeGpWdOUwxy2utliCK4B5t7oEl+Uyya8ama6nxvXtS+AlrddqaZ5nNbW2qxoMlDWnW3z68QNpfh
BjFWTWxpM+WREGaKKPIB+PC2kCiV/JM3yGPj94gSirFh3qy+QXZ49WM9mw9PUFvcgRw5npHbrR8W
w4GmolkYb1piRI56H9abS4MwM893X7YT9sZLIgPbnfpoWIs57Je2MvA1FmobcrzR4fnC1R5JP9TB
qdSvf+v8kTyjQn6s1iPCqdWS6Ug+9jzd7iiH4m/nKrxKN6II7IBSxEClZnPx21aO7Ab+WFQr+l8R
mYFEUjMgynEvTlSUGJTgfFZCtPvFufmK5KNClQDHiYcdib2ugINDlQAUC2wt6pM+I9ul+NDvksOH
OTIGVkEeQhS3r6GTIabQ2N7B3yM7uPRzgK+ep2HhpvigLuivCZa3uKf1ZGRnmFakDJH5jOsm4Wty
aScqwqWSak7FAqW6qF98R78CMeVCPYgSuXoQwZ5VfKRcVRkHuEHbTfSVYATao652F+WBKcR3RwkD
QD5zaEx3pcOg0qy1kuya0EpuR+pCZldVNrP65kGxlRGZtzIOuJyEOeUa5RFDzRpP3W1YI9/dck0W
gKydoZLIl/YHgtN/htnCs0ojMbCwLzp3hCeIHlI9InOOW51Wf8Y4L8v1xWkjHwj4jkYfiN6SX1NJ
eggeNgD/z9q/Q0mcFFYDkzSUFjIJq6lBNZeZAc+5JpZsznffSiQyaHmcgQVlAenUNVrgRGonKrqK
BcYfZ84hKhgoDmSUMmylCgFoXgfyNAe2lmRdLS4tOw12XK4HxrwwRopy0QqKVr2TDsSLxUczvoGI
X6BecHsTVeDMyAbvI8RQ36AF/s4cqmiHXbsQZWMc4kPoQypkV10K8p6DTlAQBQsibxZz0o1n+1ak
YBRRYYFQVvESnjK85bzcDC/KfLIL/TUeNzw/Ws8GUHt+xVOm1fTR7l5SvD6diwAsDNYfHv5RqbIX
x1Yu4QlitsHxwMI/1aZNM1WZMUIcPZteX8K/njM4pvi8k5ZvDkFfvf7Q64vnXpN9K0YHzJdIN2Ue
c42PzZA9FKCIJL9w8N8x1QGqZipD3kW6ZaTxnhtyqnpXmF8j6l0hsKXJJAZUC2axds81KWVO0UQO
cWkTXRjUg5X0gxXHylea70q+yXrOnTjXgVz8EwVtet1GIqLvWp0CsbB+nPQZ9NJDjekmC8IZlKkH
+PRElHaTsWGQE7zNNGLKikGVN/ICLVsapU7l5YU2reN2zAupobd4uO3r/x6ZEan35BGZLQqUGwYa
RYIBAKfqtncWgQa2c2XNwMwQV/WHY6IsDfRncUqfMWMRhyaiHXBcKxe9jv0D2ff1mlI/JC2ald5B
Yv4W8Kdq5l7TJwwts7AAc/8In4OG6fMxom7YegS8grLhIH76ZZO9m6bQi69laoXhKVGA2NTxbeZe
dtIKcZbRcNYAOONlnDa94wXmCe1alKtM40IegaQTL4NZoPV4bGEJiWVSherqRn4BFr52QEwMjBQs
w5B+IiMf+ZZF+6IZRFFAxX+O1kHVFSDTuh/5GzwutMHmTK0ip94zYCTs90B9FGlzEdnKM/pHTRHX
wilZNPQuU/DVwIxHy0wTIJGxlp+9sdejHasDflZAKEQ+G4gTEBKMJe95Y/TzmMZbr14Uosg31YY6
KtPnd/sYhUtlIo7iquSS2c2xuOaxnQONsQJHY93z/gsgKWVjtQ8pJzazew3L5GL8wkiL3YsuVeCs
NZ/APMs3dm/qhFqwGB+xThuDpKQSM71LdmuA/tXCn/PoungmZf8EmBbQKAyLOaKWaRWRyAomvAnw
QMsEybzInEA7vA9gRG3p5QgntAXWxtEBQFGJs9dmc9r6Gh8xBcV+qlP/cSHUj6I2fseAEdyGYeMO
DIBg/G+wy4WwBiAjBEMf5yv+x3wQU6fiK3MALLgHpU7UdO5HZ4dXriz/lIClE4SKRQroH2rvmf5M
iRMyyRpf46R+/9BHt60nlsvri8zFNZUPSizUF6zuUXkaTJXxLD+NcvQ2FzbMb8L2Ed7MlIsioCtO
pWGTRT3b7RBMiNUveUkDhQLUHm3kqK27QdA63NkHASp5rX2QUpXIa/MOAL4u6GQ4O35aGR6I95zM
7OS6lBWHGjejn83N7AYL2GFtXvZ1vEtLAmxRBOPTHaB9e0QWcje+GLeHqxXtrHIDRGKv8GHi0R4N
VYeB+oLgFJeZF7+4pUw5Me0FbjEDPLJKWKQzu0n7Ib/FreWsdCKP8wBfDJGWZx68LZ3Fi/wQ1vEA
3ATI9HsU63qwYfAJ2l/ZbyjujKtueAS1DeGpFeayB/cu8wKMP6YFLxvjsI9Qwhki2E2RWzWVuXrr
8XQmm4CUQytFg4/o7VqP4yZnxc7sdChQ3WgYKyC0rA4aV9n7FboXZUNQVs7MPQEcR/bwhKJ3QqQo
G6Ma6RxYpVmXSzWpj5rMuTQ+07oo52ljZO7sVA1oByC/qoUa1eGUk4xJ+hwrWWaK8cNFkBGgQ+oL
wn6ZMh0RBsvMwg4j+u+/vxuO6dFENy6lVg1W5agaahlt/7Er1iu+p+BQj5rvz7Dym5HQPf00SeUX
wtBOq4l3qIGGMpkrgPwiGjvJYM2HW5EUsKZaeJ8i2q1aFggsqjrSqRumAjDCSZ6oaWaSsYT0FL8r
yfd0oUzu1VkpKGQqDfx0MAaUN7xTxtfdY4zxA4bkdm3ydk1K68GtQQHj8izTwsGQGhruQbnsKQDP
ThAJ4nD7U6XgdSmmtesRrlgPnJfDz4Hd3Q9dsK32Kuv1EkVpNJzhjmBjQil/BRZJa7VAWDzkP/xB
b3AFfvCPH3CxCQ7TmycfnxQaL9/YKjwinmSpIExMr5jTQu48nTfccLN8dIaobH05zviO20iRAgW0
kBuPcCfkcUdKKDc22m3X3khjDD5I8odfJOYBh5/vTwO5yo2N7d/balnvGR8wlVa1H+iBzofqCLKe
IlN9RZTKIAAHwf7g52NQO7G/+id2NmkeAS/bnZPwXKcLFlnU1SSFUKa5FnY+ZO04WXDIRJlSvcaT
CdAi6sATEugLj955iKB521iBRln6GjF6+9+abX09CmySXqFqafCoQEDYAIFQKP5k3HYMZXqIgxFe
EEXiKU+BERZeo2JeeB9T7lTn05sti6IdhVP5zNbgSPj9bC35ZTS2GALGBb4VcHMDrI8gV8SZQPB8
NE2rAYbWndSARvk0YIJffC5+oCpeC9PdIs4T8Q+//1a2/OmaBwNEqB+4AlSGcyzc8fzP4isS1KqO
Qklf0lB9ACtccHT2AqdPuw4I+qZw6rNMt3flAKD3c1RyzcW9pDekmgb0781uPATBzBx5nd93dcpM
1rYXoeACdkdznzPGq84pufJc7rtW5T2LHaH2EMQf6tfJiL30596R3Y3x63tTjHTWrczaTWnCPOWW
gwVAYPBtpWZvFEapYpqQGJ8rtBF7gVEnpdzI+u0IsW0640LcCcec0xan9hNJG4PxqbhOR3Y6gNrK
xBq/XxCZKJTcD2vEGDJxp09D+GiKywFXJQTni1TgrgE+izYvD1L7MA9WpqTjiKBwqZbSF3HOT6ZG
LBCDUhtQoStp1yusK3ogAFm4UxB4maHGNvGRYEis0BGVUqrOflK5eK7vv8g4OPfBKkKn2JYSJB0m
+89zkMn6qjudrq9m4GZCCB7zKaNfsEmE2q6PT8Mm+mufWvxi9AcuVlO0YSXem93Of+G4SVbgfu6B
/e2vO0/bIiyNEMNYLr/47jn7C5uX295i87mMz2ODwpxpwYqA4wnNiLkGDOekpsjql2Cy93uFWyc7
NQfn3Gya6iLJFQPJpW2WLbVNEbk9Ec4SCllj9DQRDkDiUVWC6wWAvY7JXNlBLegvZ9uycMH9M4IW
AojF4P8VKLLB3NqFp0OcKiUy+bHTB8Oy7iaC1dgX0ZqKkCIn9KDnrQClZ/+8UnJb9TQON1f8OABN
NFcbEaosiG0DJb+JFiNr3iE1xjV5J1fkzVWQzA9RteKAgz4yid5vG6TG2NRECt4EayxCgUrpoKbc
RbxQNnGPcjCAUMBfP0MiNFPflZ7jjQV46P0f1Sg8XbyahAiQN39PkY/rrRv1KRENkaPTdA/cqC4T
vn38Z/GlCW1SmdpRE/l8uT5RrxDCls4zONFFsOjqd5NmwVkcLDMakXvz06kcVPITnh4R4ajuSIrd
SVVo3vUEeMgL2css12gicL/jtP+iOKhTnrzce+PUnFRWZpNq2g+3fV76hvCV3Mt4nqTADvu19LIX
9EjGzzjqZYRyJ3ngD+/ExdLPb32817hcH2DVbIYnjTfX6iVaolDdczMJjc6pTnnbCXYDXC2K0kb0
SUvn7qOdEyNW10ttzH+x6ThJLk1Q6FfuxyK78B2O1reKkappRNCCNArayltgvTgdKLU8JNP0x7Nl
P6/yiZtxg3xANrL1zG7xcKw8Y5qk7X6KFUXQ8buawO2to/M3VTg9bwYW60PKBx9lEnSNc9wN55Fg
rfxiCG1PeGKvn4Ahv2cAKL+TplAhLIJk1Heq6ts63GDJr9p0RzpV28QBkW0pSL6D18rO/NULqPGT
+N8L6L7J29Hv8xCpGcmpRV8u+XRweK6VKFrNIDi3M0QmVS8k/uOelnlwhzRy84nP2DYGR3kBfgSt
djB0oJ4Pwem5N5t/qiNNV46k/n6I6mFY9maKKVjRm4AFuOqPLTUQs6Pjt0VfZkRyX3AvX95mrbQC
bAukThZ71fXP71dlOZJaBANpYDL503OFfGLGVA85kYFLKvkXM8XvJeK3kHbE0W/QEVkqoEPg71zp
1PCRniTtahJ5V8fsLJ0/0i0nnd+HoOuEjmB4kyue2bhZtsao7eaqTMng3ImA6QRKp65BdSREoKut
7xekYw4FArq11t7rG80piZKOHmH577GNfgY3/b01NR1rj2aACGguxFlm4Vhq3lmFsaKRA1foTuPp
jbR1OWl/ncFWSr2D3AkiQRLb0mKHhw8WLhVnHGd96i0BpBZH/a4NZJhoVHgLzDSJmsjtk2WxQTer
nxxemgOKBQ4BKUs8/QKrusKbqwEy6rgCskj9I3wqyMeptmQs5rj+gP1YFqfhO7ggzXxUE8vIbBOz
STfl+FsPQY5evny74rhHeOiSViZNEI+u14x6gYENAWutZxWUKdSPq+rvetRE5TwtZLXizbtIXReq
FwsnFv4AawSjzEhgB67OGAEjRJ3Uwht7EwcY9DFe9dyK6xTtYSeMQaPDVGoS7102uqQ68g89zxkZ
VsxKwCEzJvaQ9kDlKoazVUlyi8l9M2mWyBsFQubbflOqOhpGRHKZxqSsf1YUZV1g+tSITc7/I0b+
tgntLAJ/QxhphA5U8c/gr9L72LlDBSybXQ3B/DKfeOuKGxEY4GjiRnvVMxSeP1qHgL2FTOdvF27V
ZROUX+crGTefpAo2jF/1K4uKsDjkuym9fcIgFEV3ZYZQQy6ow/rtMPyV8I1K6dyN1a23bnpDQxqm
nQAsFWey/fx9Vu6JTMnEzeZXWTJtmEiOm3RRAbNGOSt2GXhQLoWGyudU1rZ5Cu3h2UnxjHJk908H
AsawBPLhXTe/bBpgx+YqsjTnsMcDQD80Y3Jl8iN8DV1O+/b5Uq6Q7EV5ZIwNQQqeKUjFTaJD3y6O
81nXyEn8+KQO2y+E01KiuxAXzA3VhAmHBBkXtrQtKjCN1I8b+zFNyg7C1RCEw1ivIrW0wzWz3H82
JcnRnC6Ncg3vFO55gAWRTkLumfbaRd6HFMqw3uvK3DQ1x64DFQFRnDf8OvUxrwNJWqHK3I3xpabH
poApSoC5zYMCb5qmlxSYtlIOFQC75a6htoIjkL2cQVe3zk9n6Bhnw+f15i5+gG0W22Ko/UfJn9ji
K8MU+mLjzeQ7Y08eEFd6vm21HCbzEDaKfYsJnmS/WSmCOlHNkR7yj4JNA1rWnJS1AL5NoGBPJ5Jn
AqJot8khVVhInkxtfcNj72TMeOyhfanUZo5T5IzxjvpBzK3mKHqmP5lTlto3/keMp14bZaiidkWv
2VYCYraMmhju8BLI2cTPbzj0lYJpp3yK7b/J+6fhIXGYFqH4I1SoG7z0hyF7uhK1peYKPphCwYQ/
u/bZmAd4gRN7Uu6oAdIkx47M+V2fDOg11yenNizD2HFXqEYhxem1D2AxXlfFFmlSo0ISPJzSrj0H
M8mc8rXPZx0LJZ/oz1rNPBm6PcK0yI12TruRAz++ZOhZi553ON8LSkkBfgZ0iw0HeInJbuvb8vAM
sPJ33C75UDCGhCYNz2OLOXuU+xCz3OkhZLrdOddmTNXYlR2CUFCKhFge4Xz6/UyRjtaSSMaGe8Ec
jAkZBil0AqGSnk2Iq9FmtOXC/AgzkxXVwmhryMLn2GL07JA36TuVKpB1QE0JE+OeghFHJixoh893
seedsxxQjXyXFUfhVqFM/FXzsN7h5ZV49Qg8ckAokM9yiwbLQqhwmzospDBCPwcSlrdWqXCE8+F1
0i6p7kyOeqANuPZP1L0oqk8tKW7b7PCxadkYf++uB5NQ7Hgnkh+aV9cZdYtDhMpML7sa9v3OXLlY
dGwJJCIgswTsyeeJrfbYJHF9G4d/Va0+fcyXF2Ertb9LEWKqDODaBUbd25xNstpHB4yiKasaaSAW
Aw+ZH+DyR/Ov+6L7BLKsYuncFashrPknsi5q4M1o8er1UO326ktfVrE7Sd/uBhdeYaipvIze80nH
0nAPuTXUmI4mxQy7Q/JE/czqaKhlGpC6wpfAmA/S8KCndTi78OypNVrycD0sDPfyVHxpvLjdgSQS
C8QhAeohv4Wh2jDhPVd3lTPshB1A1lzTrjBfxSAAXrHgw7ZyztubF0EnoPo+i19FfbDat/7zk138
cGo1IgNtcQ4WcDRKzBQxDimMYjmCgZDp4853U94At6YWgNrtWGu8Clx4iYUTWeH4LQiaxC0ia5A6
x+p6t108GizNoTxUysgyVoFBVihAkBXaWtHC8/jRZUjxGev+Bx7TtrofEmxRDFqYPz8/tJf1Ex8f
4qSJQMNVJwkcyPa67S0zqGqZEVrJT75X4lA4CwP/Z/lCRAEs7dP0iXJf42bzxogioaol3Wa7z9Rq
APdNaj3OML1XSvDyvA9So4SievsICdE12wZfWdzkkQa5OT4sM8FoebRECnxsGVYZ37epgTo58kO4
86gGoeUQhaacqgm3QqdGvJmCvy32s66Z7E5aWkxwxYFHth7szElOz/84sAqSX59mYSgtPR0f0E+D
I7k40ceeOhqIHPgW9Ii75syeklLodN2GlHbf9Nqj8qZHNQ5logsPeF5eDZ5pd+da3XL/cDRpXqlc
AnpXjGRb9ZsqtIHdIL0VkswnqJp0AfQMiL8gEJGti06cHDQrN33YzjFOHThlEOH7UnjAsJ+pbzwO
kRhRKcB2Q+UNsI6AWlz2lSCwY+89T4Bnnj28DHCl6sZbyYzs5GmG7nXNZcrQYL4y4hJ3tm2m/yyq
IgL6nnaIvpO3rAHk/DXkdLyEDjMeMBhJdyJo+PCGmXgLEXkPOyYsxrn1ls1OMXrQ2UDq6pmqaCgS
5IvRpJkfaUUlMUd0MMnHBt7lzKoW3EhpOjXp2mJsYfx9DarciNYKuKat5v2zYhfFYdfljCPh660h
HD0g1knyhLEbpc1Hb0HVq1TAs5OlR+lwFnkc9prQ2saBiz9wVsbeeTm2UXZVuzkjkrHKMCEZcZua
WcQ3ajl681J1C9jqtva0r6tHt8OadkAGs4FrtjLVEfpAFBKdRPhfANZzFNEwq3LM/mx6ADWjUHps
/pQsJqPUl8O9hDIVxsVXdKT9WCL/uG+K3VLaQzQ4CD3AEcDccQ+v6ACn9Sjv5yxkj9/pxjbeQbVy
cFBOv44Ne1Jx+rZvzayqA7HtON85od7crEOFRN0fssNYzv2REoV4hlpBRG1DFkolixpOR5rmrNWJ
ZhkRB0OKO6535cXypNgEvj1DQdLYTGHdww559o9NQlKciApaA1u0Wywuu3GNZlxQMB6PHicOONm2
R2J7241YS8zLlPTDwv7Yy3Blk2HbJ65C6wdROQSbNwHGb/7eAsEipqpz6ISTXpqtEQTx+roxcQ8B
KDrCeyNUbi0D/t5jigP/2U9BbvrgcG+2Xu8TzWWCm9FL5Ib6t7kT2lepClX1JcN/Ujg6UqWNR4Qr
hnnzQzVaQEY2gcMxN4oMrF0Dhv3V4As2LS3TwfgSeompzIONZ7PpK0DAR9VqnbdKCHV/8cWXmwou
ZfJQB19303zG5mkEjsJoyvpW7DeiBznX9WfkEAwtC+KmYaiMyRsT9y/3aUSQceEwbzpBj9Ib5HdO
EgX1ckQKt0U58HDgSaIVqm6orIv/+CIvrwi9H/j8Dh1ns0AxXXz1KFsyFVA+m+YpodQhxdrM76q6
H/ER1wHrNwwyU8yj7EFBwMTPfqQuVa75wVNTY2JwWBNSmningg/Oy2Kc0VL4K9d3B7ojwxfzcaBE
GFSpTohn5R4tM36z9VUrVf3RKkExd3g7YI30N6G9D/0UfJ3DTfsjgrSu5nJKdateiICBPtkpm37i
FqI6zYbmOrqW++042H+EazK1xuk4xJOR0V5ViaoRx/BanHzscejziJyZ1BSSQGJKPKke6MZen1a2
Hl1B3X++r4kMHTNAIWuW/PgjIZxOeOaFXURwC0HNAdtXe7JGDQf8iiM9BmDZdwKun5O7FcGqSvn3
pwJb3NRrd5x7ENVj1UoeodoDPLYKSFQ+uFj9ZK+7qFUeJAVrd6sN1YZw2FIbwRJCK1mLRRKGud1p
5mpZ1smYZZOIkfVztWQECq+C9IQhaO/tAFnKe33o8YD6w3FLzNM487/xFycm36kJTcUFIOUF2uw0
iWSPIfLoTz6V+XuF6o7rpGvAALyi4ZQNU9/Nzf+WMstvEqS7E+WDFVCpStPpttqX/x44wQbj0OZj
OA/rDd8sQN+Bo42nlH4qZnjP1l+uXOaXrj+6AR7xW+gmEVUZ2ZqHIv7g8LMxiUnXstjslQWfDECk
I44Z1O6VggMXmUndjCgZ8VvDU1r9PruMfh/8OkWpWrZTu8CVgNYlBgzBgwZErI4Y06AKWsey5nh5
dVLVVBfQ9yREPUlDHySr0Cg6rH/NVyUs6CvXogXj3OOEMMxcGQouDFmYunp2WEQDbFKC3D25B6Ns
2J433OLk7guT1Zq1lLAb63SC5q4IFZ/tYndnGyxWOkiSOWahzSN11dunCly5LIafFKpTe9SqoHig
d2ALT2d+jqUHJh0r0ij7FuK3ciQ5SgMj+yWeEjGwfrmqSvuBkF6m++TDTJDC0IdHgAT8Je+6unir
CvmbZxr7gWJCLVIQ7i5WM73GAH5yR8Qa3z/S1wE2KF8Mrr19EXcw4wcQ3A8aIy3HecesvJvrpJJL
8WaN3cYO03YnD6vegYA0gZRPcyLpqz7kWODhNBsWLhvYmA7Hsm1i5jZ8tPLdHudt7BkPU+CbYjsj
gKFOoEhqHkjIegv/EJDRaI3uhPb27rdAtr1Y2yZeyXPNzbkkctujTpaok6b++L3FKiZiQrWQrjC4
tTT+vBEcBZKQNdBojyLxzcaktklGnJlo9v0UGdW3Ku48PrifIAS/ZbqzwgOKlUnu710Uyjwr0SON
UEqx8r1dG8sPiYiCBeoFs+MpackfcFxawXGyVryPHLchwj3ksIzwJkanxAZb+MoF0hvrpWGwgGfj
CM3MhrZ/TJVD+0CnFh+fTxB3z9RvoJ1zIPfs3QgI8gJSGiMrZ5CoovQF/Isvu8zx+KMLN3z/kQwy
ywyoTmY4YGFfOM7CPBkcBlF6YELNvnCi2vb/uYhyMTyGS9+J436w/1Q+4oDiLHFcmA8Usw5qYCOE
JyO+32CYoTYaahQ9/rV/1OCRQoKJJgg+ViUA9ETvvwGRbtvZhyDQe+2pfpQUIHl67cwVcMjPLdfy
kiXVwo8zg5FEKhteCyVl/pEvGgortJJuxQfDdpPKQNCciZOES4Z06lRKhinixRLlEIIV74k8xC3h
kf2LN/DhnpjshXzj0jF327Rc9CJ79PbjjoflOGx3y9c3d0Thsrzg6FjVZYM3Kl3Fv19EsEgBBUYq
lau37JqDh3HuNjwSfjtgdHEzQa4l7acLgZxT6DKW0VUKVaul6w8RBnU26vYSLEEGxNRwbmVHZ8Mr
t0eQhNt6yk7hBf3OY+WNnkzuzg37gTSs2QfOMICVhsagVsCaFmrBQ3UJDJdVarcsk+xCMJWYZp+V
yE8VAg5doIpvuBHEzEuoCpDuK/9VCCc6bVa5vJyjyKTkFBRn0LjiGuz+2Qs5mPbtDWuUBys3RlHn
vp47kVWn0Hz2bRI0m+NK7E9g9W3ztFmzUeVa/UgjnSkpVP/QDerMYgsaslbozNHB+09d9hAkHVkC
Y+gBxCds/8eEwudTPBmmgKKQSR4desQQ4Ozw0dBRxpONFizXu4wdmZhzUjEVxpvbEGkDJ1avHWLE
eN+47caCkFB+yEElEadHabJUSo1CxI1u4xM4ttIzeFhRHAfHOC6LLg1bBr4EnjCsWtc1K0caYxtG
/f2wI2PhpwFUCyASiR3nDa9RVjMEH9LAzaC/w9DKfxXw6zgEES7USOqyOnmoh+kuMW/VuYrf3A3r
DhBBx2qC3PR2oAssO8yQpeuhg9AHimKdG4obQy4jLWUW5A/L04tmIx33NdNYfv+589wqTK2Vaask
ItiwlsT4Li1+PGstRvdHz9/tW3MU0aiQFzmbi57k9R3BgexeHN65WAmzEXq8X6G9k76nHz04iFf2
og+Ftuhb7HWHaL0lxznmaQ6C/acj9WZ/R/t3hNpcucZDHoWsDlwd+UdgZvPV7W7ezZiFQ4ttWgNt
a2eMsX1fisJ0R1MHXOfDVGumXdY/QTHVHOs0SluXzrY042HEN668mUKXWV3yA3UH23mW6bLSp2eZ
x4QwX4OqT+CdIAo5T5YVJt9j32iRPhRTdPalGYTM4VARxnagxdpoemjGSik2ljnqt4o18HdtXYja
fGiCXhUO9hJ3Vwuv3c3letKBcNFZH7rLkcvwkUwDssiee54drHL5JvcfdKAs77+c0mhHPyA1ekEo
DccS7b93vjJrJKSv0OrT6MhqgfMCha/cKv1l065h7FRbUHrtRBkqxiY9C62Q/s2zMqK2twghX3gr
FNB3hAmWUTywaVBZvU77XivLEDFa3+i8JY3IUYkLoXW3oxThR4vKvozv4PQq4i5k0HznRxgv1zrw
UWtuQAm/Na155D3tl+8+vQMWHoJUWSK8aTSUPUIeKvUKa0Y/hKbvukfIusGLpuolZ2l1pYmDNsYC
Iup5z4zy4IPbCqMAD0XplpF6Dq+0j8DMpWVR7aXxl1Ywinab7o7d/S1HKnCouN85P0nNRzaIchJK
BUC5JG0xR3T1T0jRKcJgwN2Q2oeYYInzJ/O9ZOPBj7PuRsymZiRadO2XOfbnWaiqwzBNjtpbpzHY
TG4FyTohgO7AjZOCuNne0PCzz/n44JoZX/TFizwI1jbu5qLl9P46gQQn5BUkx6E/vwxki9SujUwd
we6hStrf+qgEPmCbelhToiCKzLyA/LYPswGZfLsuk/GsP7waKAi82vOddR0aIWklqLS0a5PXn9Ki
WKNNtY6Eyjm2X1vhrMY6rhSJ9sekkmg92y4T+yfX8NnjuZ+f/2kV9WhHY23hP1pn3kea2JAvbeGT
Ntb4md2fHV2t2PGy94H2U9VoKHvhljwwaGEcI42sHT1DdP+EJsQy8CFa7joNZiBhPj5OH9g7dQTQ
WdkdZ8UexcbRQObkkGVp/5pUNQIbpoL7d/ZIPSgOeEcdeF1PGomuDm9ewav3WeGryz6rFZRlH5bo
nYtwmMdyzmw6kNBVeDhSrnJEpMTnJm2M2dIv2qu2v75tVMPpdxP8vrUfIpbnpPdT2A8Rp0CcUR6r
rywKEkzpw0q3YAdWJAUHd/0yYp6SZMKk0jkjtdf/rXiowPhe2KEmV9ME6DNuKxxCZuJojpibT1lD
EYs8hZKyY80Zi6l6hA1BqwwnSfBKFov43m+gAharDpsJrgCLyddWfs4YhfsFRPhnIAIFfoLdUvq6
QDtQgtnJE4bixkVEi73mRGJjM4PxsRp7ZIPpbVdMGhPWCp8LoFXXXAtncFVbk2xQkCLwP0DnHRQs
sEs5bbGHF/hXHplklBxzCtYpRxWMlUGgUO3Cv1kBAli+iKta4zNpucY0d2e/4esVt9Fdayr8Gia6
j6btwmERvFRJp/71U/AjCf0jvFSsiHUX0Yz+T2ll8jkm2cFiypZkLNNOUs6ZF/R4zSOfTgEHqD8G
1iW+0Su+CIbEoE6VQ5Mq0UOphv5ZWxxx4noyIrEEHdvxVMbx5VNR2qYTAhPqBEZetfSTWc5cB5qn
5ITaVzeOikCEBlWDv0YhxayQcL7/U8fM8SPunQTbAcNXR1IkR9mKkx5OQFumQJDm2c9Pc4JbZcl/
MBf3fVibVmJ/ENnHl7sGRfcxEcgLQKrIySJMC1HrccZ9ZxfMicMuFcuMKNuJmsIr0DfelOwid7Ke
zW/6d8C2yItOEntlOE6hfXNK0DRsuCFTyXtOI1Bp6thoAvBFAp0aGbixvwBIjFgoRhhHT4SI7qad
s/FU4SSdaWs0+zS+hRwXEGL/Ey0kYqG8ZBfoU12Ro45sXWcqBQ0xWBb8VTCEoT9i5arGofpTdYAj
SwrMZRaf2JzMYXzdj6RBl1e7wGOekTjSObBH5Rkec8ABQicOAAMfVcpP0nkmvCnxA0lCH9rfQ1yK
CX64QE9xhFp8dLaWBKdrgvmTsNRqDx8kPhoxYx25iO5dARlpxlyl4U577JIphM3Tx7IVGQ7OFZTU
m+qrSsvInn+9tqKTAUsSQLnmmBRkzfdCp90vgy9ZBrYDezLmOOT1LoEqrN883eKJ5A/68OfOM7hG
a+ey4YlJM6NJl9oEq9BlBXvGABwlTXBKVEPYwFNx58RhNtHgf1SJpgYCAd60PPGJEXZj7Vw2D5Qr
Sdaq8z/GE6RUCRntfcFqI4r6asNnKZShvl5F0NnrgeJk+InYIUpb158UJEWAqA/TLm7T6O9LiT27
/2lXhM1J6P87OHv71+aqKWXcK83DHYXE31dkR9FY3WCsBQPVLIpqxUvinHA2N+GxpjKDnRag31DR
4ymgKJrf/2evz6nicwkLeAqbltKciCg4HAIn55y7vCrAZ1q++SYcCJf2ZGfZ51vVFA+HcYSoLbT4
y8QVPm2xcpgsN6W0w0YbrtqRt+je+qpooq6wZGAo/94no/GKWam0KvyUGWBqlK+4pj5/yonWJCWS
HjTmEprVapM+34869eQ56zQn6aKILLm3J3PhTJvlZOwUqDlToC1tmSeRSSy46O2jqycGbC7+3H4v
4KuusENSrMY7J7RQo7e3gcwTPWobETJYBXNMmXagZRUv3v6zgon5ZYcafrCD/qDT+4YLDuSQPf2/
ht7u00F3uyS7948D/fmO6UGmymoeg5Vk9D0TVDCGdyDhI7876vfHtqOwdB8Tj+EOvIplOFpFiWhN
wUy1USdhHxD7sKVNT1ruv314QoZrQweqRv+weonmfVmJ1MwpO2RPs6407tsptzOjHFP0bNtXkay0
V5m4uquoKXRqSC5Hm6pKqFUcZeaazur8ATQoPQ3ztM0Oe+bUDV95+VZ/k5UdLSfSzHOUkA00NhEu
yR503HKpUBte4EopF60nAFfbG4SmQc6VfRoC/3EbThYVwZJe+VvfiIuqHH25LlN6JsyyvM1GELWo
pt44gSSdr5D4mcfA1o5BAvjsBnSsI43UE68idksGrN8kizbwpKMumMshj3711xl4Kp8V0CFe3+Ou
iqzOjDxPe1jaQGvoeb88xs8P120l7DwxFQRRNEMJoqXhdQxr8tjbrhw8RyQZUB+LVtweUX42kNfK
3EXe9HYcClBue/9fYvNHHrBU12x4EaX7sERVLRqcVqj1bR2QB4+KUdK1u0IgdRJSb8aVPtiTkdmU
L4DkSniiHp0Ig0SkO7bQbfiJ0YqkFNqxvbzJSU1Ed7KFKED5FEnxAM8UJDQE2e05ErNWU4kM0OO0
KSOR7oHy+P5+eyttn1dK2DX6OfP9gp50cVYSHzCIlCXJ0tKppIFzyQXTjqjKGrfWvWn4byHjgsnF
vO97KUbP2MaQVPu8faQ8dKxUAYnx5Kgkbm163uPMoZ86M7cT1QikRJUD7l1laVLvHmQkcdeBdcr/
jUm8hN+w8V9KvoGgk42+LoRnaQzgK6Skxgp49Cgp71pWlquN1qSlXFcXaOmp6fvAlblyWMZZlaFZ
g0j1T3tNBzKXtOI+xQd/zSNqXB394PEtYvZbTRgjIEO8O+wzOksCqOoZY+TULgcyk2e44KXmNDFF
mSWXn4V5GnmDyrmhMGyNdJcpnnnaj91wOf5UeWYWruVsPJ9RzmhDYgOLKO2GV9bA3/KtiA9tSspa
xp9955Zn1pMekdfIquw50CRu+8kG6PieEjBHurRjxyGqRgZ38BTBYoNk+tYWli1reIWKGseoaoKe
wbk11hZy/kCY4F9Er8ehq/6xrd77C/eX3jytf1OIVEvhox5pBHeB+Qz+A/6YvMrt+i1oh/GZgEBK
TzTwb1Ii1/jTLDdepOly5gTpyssZsHuOpoebKIlVJWiZSp1+IK5QsZzDzVbzhsyE02eXYOyHV+RN
szajmbOXUYJFnuXRaid81E2Jx4E8GlUwkDO8J+I59bRU2E6haIoTpm29bqfu7YiqGpXmnCAdNFJt
XsABUhfgLjU60Sk3+i+mzAAIcPp8P5aXxMyv5b6qhbRYC1pIN6dk6+eqXcCg2S257CpZVrvbvfbo
weQXn9Nri1Z+NoGcctQmF8PaAUOrx1ItQstaeujLd4Em5Up8/4x/uHVhYXd6nXvT2g11il4d65WG
KdkAvPPU0hBjZLyf2vm4c331RirN/z1nBTz1qDA10DBZ4/VVuIzCFVmHKy/X+SehL5BKfe46Bp6J
2+RqphKoBX9WrZmxd0aJ2p7S7j1ZtAWU87tDqWdBouNpgpgHvGGanUnI5wRbkt1Antzx2fwjGF+R
bxqX3O6lbcXnMgOnpiSdeWAE42jo73A0DKe29DumN9ykqMiNH3fAS33TlpqY5ccpD/xLUaYrP+Rh
w+C07o6MKBS5pnWE9VQrSR3dAyHWMov73n8zlEKJp4919ifNtAXVsfOUtYhc9X+tRxycIBYZMU3u
bHdCh1PxAZZj6F8+dfTjn1P13ZlmaXkm9gU+/44y0NtdBtcACuCZm9x55IJCMViWL52RF3EFB19c
6DzA2DFgv5CKdeyhqXPApwPmkZRnvlBq5wcYsLhtRcv0pOqTn/RIsNBsFJxge0l25RTDYEQh9Zk/
F8Wxakuqnbg4ZQVhQFEeCg2RnSoj4kU6n8aOggQswB2dvuu2mp/gLKDXyAo6pKkNuLKk3srg969v
ImU8i3KNUrm0Kyd3cdtpiWFOrH8lrYWd2a80CqJq52IYTX96QZczJY9dVHWn/x1y08i8NAwAXxgC
gqh1uBglnCaIiD810wKgBylp5dtbb8MZLVrZQ7AzDMrQJgehz8X9dhEr9/I1y3T0Z+odLHlvfIAX
P9euWY2FUoPyhfRcGXrHzvilW9X60JQTSvIJdWsD0WeKSBWXzTQme2/t0p5CVNxNKGTkZ5Q1UFt5
6+8XvUIWk2eQ3JIKMjRUMyNUUgrI/hrUiuph8VINQcInbrJ45fj+5PT0s2yUHwa8QuAiIjUUqeIr
AMDRbHxdYrzlfx5ic/nj9PuvFBQp1GSAP5S9b9GzeY+esmhkdlyk+5LLBHi/JiMSJwfitwHHBI13
GM3FWCQHjXNORi83yWJkTYugk7JVy47KACedI+QX/VzUY6ikig+O9h+FI2gOpO7CdG2REGR1G8sP
BBge66Ahq1a3S9b5T/DsrpWCZOvuBLBqpwUf8BZzoH7jEdNJu7xshm/YWOYN6+0vIwC5HfojAmv/
wHfBv0hOpQ9IDHo8gZ6s45EZ5NoLdoFHnaBC5VoE3g+CYUUqjBVZWuUf3mcRho5ik4QnsVssuy7A
xTWj1uz+QTuFoMKmIGPX38mmWjpoFNoshiGIDn5RMWMFYFFiVK+zhU+67ZjNgswg6klxDi6C3tKv
/WuDEdK+R6+A9Z+ucbTuFQKUSqjneo78Q4nBvOjE2FWxfCQM/2xjKGnBRPQ98OPZmZHZl9HUSZfj
vyAUMetsv6fkBKJwxQzy6RAKSJ/DrNsyZ/wmyQprBMXwiQZPKEfyGfITzA9U6fZ1DCT3b4LdxWCm
7mvIKjsPn3yU7baFVWNwOoFWrCanMWbhe917f+eiBx+nDwM2gv/wxMVyET5eG4L6HvCsKoU2cvaO
9jgwnezuVpSUWTl66dYLvo+gz2moXLNQO9rhmuAvDiRMGzkhrI9pwXtKgeJC6KVtcitPls7yRi4Z
E41A75b0mf+62wVGeKr5QVX2mWJwaaw=
`pragma protect end_protected
