// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0.1
// ALTERA_TIMESTAMP:Thu Jun  4 11:11:14 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bTm4xOPpmQcWpYnUSZ9ZdN/g1ZbCZSOuUK+uvyOxSIwcQcQvh0ib9gQKH3ms5Kdy
Z8I1z9XpHrOVVTvUxZNYpyaVPQHOkHGWs4Pm9B9B7PsRtWa9t2JwrJ/54DY35ctd
kJaSLq11r2fn17u98CIivi6ZMqHEw2NbtxXDfhhlO6M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11456)
vlLGrej2AK+tallWyMGTizljreW8SoU5FhHAhZmDQJuPr0747jS9Xtsx4nvuODOq
iYEhvNOVTB9+NEWTJzNS24j3cIXpTSJpNvjz1k0DCR1PHsjTBF2K9zWJleskcAhx
YgyU/0WnTkfy2Zzmb5INnDj5o0+U3Rkn1FxFZheSjCPIfTjq/XC0xPBBzHvPZVaS
YEtJpCAtMLpOmNVMXGvqgVTB9G7Xi9rPEFvgHe/+zTiESzU0Nwi2Cx3Y0dmnMg4I
5CSwWfA7bNkYHYGlqVpADGTcHCC8cnucvGGRKEjHj9fXukgxa+lJmuP9oHS3Khwd
KsdWzOnF6+wqj78L28iqVpe6cZ1u8QxO+wCq6in9gdTLPb4baxyxW5vq8K7WGJph
fxaGSmBUzWrQQQ3E7NQIPu1S0ogOXAnWDmijJVRJ++sdC4+ipSLN6HdqUj/VRwi0
9vIWsn1mtqltNfC7svcHV3DHz3I44uQhXOuLFDTndtxyKnRLtRwOyWPhNsxm8h8Z
sEIhLBu7uT4XQZufsEuuUn56ZFYtAWNxunRoX2z1ug2ARj8U7d9yiv+YGx9KANpG
OMsfBQiVijM7+655RVKwFmqaMbRIlGisJ4Hz/Pk2aOvB7oigp3U59U0kA7VNBd8r
rAzUWgixgk7MuJFxRoG0wRhWAa0XgQJwlLk82a3JlR1uMtofbetZqmN23CnOUCoi
wXdqC84rdFsr1si85a9DxkpM8KQYxhPPXulFMhL+abf5QsZZQTdZEgosyonV9tcj
r4zfy9pBgJ2dYigMb29IIt9BQheooKbgm737FTfAiroYFo4HGkBg61Vr94c92L8E
mtYNXh8EqNWlESxPYO3Bw839DNXOcTnlV4dPStbySVWwz2wUwPpKMuYSSeT6FyLJ
z0q4CcEMZ6bd5XKXDooqFguz/TmvvdOWYD4d2uXzawInzUNGqBuFmyO/C0Q/JjKN
dQH7HIwQoI/02d9Y0ZhFpIAinkIFVZVwPmQgL3knF01cMQsfwP8TfnQLI7QFNDpE
7T/Jtagsn6iilJimIZN7c5xjfEY9CPqfMt4BGSDyXRX/SKHJ7CJHLXX6qdeBN3QK
ueUZc4IJQ8HI9a1NMZPuEkuByVSsE6TZ7GL4WwYKb2BiPYArf8jc1z5/2AtNCnqa
J+rwGeNgh5cMhuKxP+x+WRzsqu/t+3zkI3H8vCcv06iJ3QrushJg7cy0pUMRMkyM
ydbAITJDXSCs1yCiDNco3j9VUCR4gWCwmBO0CVCftjrE1rPPuvu3iZmJ4DGtdRpI
UQcg47r7p0FXD9BbTwWmnKrUWLvRxSFZiRAEslg43tPcZunASzMm4ICF12++GhIv
XzGe0zrLPnlEQB15iOsd2I9cEQvEQdR3+XTlncj/01FxUJ3NC/c3//wzvGBEEOjK
ldlAzz1w27fIb51YEjHDy9Eo05IpvQjQtOa32yV8xiRGh4dNNIsHL7VrQpq1SKH4
DUgS2Ai9ovluZZO9LgBy+BcAYfZV4YiAJIMcuHMBzSKyUm/hGOpzwT9KPYljD1Sb
LQFvpDzrPEVU7IHbmRHX5wUgjVWDVKeo7CVzurWhCKOCrkPLbf1haTl4Oz4wocdp
tmNKOeJVgC6tmeHNmvsWZaiauo+HdO4ytZEhbDlEv5UdHcd1lcat6HMTzKVLqNBy
DizpXm8lQlONvUVFumCVvveriLKv09pio7oDXfd6cQ92x7GCl5nJ2d6kwfLYwAdo
qZ9buDOO3QjE5bM9jJDwHzaVkR/9ejvOHqSj/Ka49VWQaBOKstesw5bjhRtxqlMd
6u3QjmPa2g6h4TeCQfwbh9W55NclSgKe6u6RBvBk4PHOwU7BGyg5cbyAzBGLYmrk
XkRR0yXC0NjdoxrdWRHlqZm9Er4vzOOs7kiZ0GeKkmRCEx6eX7UY9rV8Aweq6JJ2
sr+eI2Y/gTUIYMe6B1ktzZNZu0jem+KRSRU9/lrrh/TxGftmILqcMS8AyJC/8xJ6
ID7Qk+DqPBLfgWy43HRF7269+YnWVwwKtpR3A0VfMTz0ilY36xTHP8f4CvF5UzAZ
RlhozlBCUVXY3ivJS9wgpBAveD7pXkJrz5eUNVEUbE7mQDW2waigyUc02pDmferO
37Wiq02xDN2N/KI7Gwp+sQW1O+RubsE6IOmhsrETQ734gsdeQ3my+yfnToxIL+tj
esXyYRuN7/qlG4SVmXfp/YsaDlt1f+iDMs5y16V7Ed9hy4r+sfVCMo8NYh3FtO/Q
Cmld3Dz9mYwKk4wOEiMLeSf86dw5zNN5fX5ytd5DY8cch4PPKFU6B3Bw6aJGbFxh
uHYFyQDqOnGC2EohzBKj1WOJ8321+QgnTP1PfPV6sFc/MpHnaiwTllxeQx8qB4B5
nuaJ070GCtg7NeS5SWH9sozZxER0Hf3+JGnelyjzDdH2w4txDYXXpHn1ukQw/Yod
sR/gC4dLF+xZ5vu6zGcp4JWl1JPN64gXNw5zcIEyHLBrNbcJgFZbK1gVv/eyIlCL
l4kaPNLvPI0WIJKtBD4DZ4vwJzllKvKicspMyuf7ZoojUQrnc/no3XwQa23bYHoJ
tfQTCq9wqwvQ0bTGuz9NMoaLj1Po9FgE75D8Xz0gX/dYCJ1ArR11Hbo1wKsp7LqH
1Bz3YJ4JR/7CDe7TAqg5/heoDW+NnWNhmfliEyCqlWnrR5cSsNoYKyqS38M3uySL
uyP1IlzUCGYOzgJD7JYjAlqfwEwXKAXNV+OGihORiRvPrZTGegfWF32hjHp6tYwc
s9HH1Mo859HtDl1h8OUg1ve0GdJD2By49yAjS/dfZ2Fh0Y00pUS7QzEZTWsn58m/
gn/YnBNSVmOFKYezgvYW27QzWJq5b4U25E1XTcK1jRc85pI37LMQGLSqxAVGCiNX
fnd5RWR2g5cfvWdC35qKJKB8DegVVUjhHnsHk/HByOoLfu678vnVdgpzTRowyHBB
Yt/eU+iy07p2j/4/IqbOlee7X/IktrkhRPHiB64iWxPXRpIIOJSWFPlMxwM0Rw+b
FJyCWeTO5fnJVrLnqsKOOEX/kHX+p8LrSQRJYgsZvVwwd8xmIdYZmJgX08RvVDgj
VoPvRXFo7nWP/khI1Kcndf1j5wFwDr1DR5EiNC4UBfx58BiyRzECHw6Zk4l12Jts
HOePcZGFVCowP0SCDDv/kHcLZ1sb5i5xH0KJ7xu3ghyoSu92wxv3ZnDSU1Qqxqky
tSCbdGvWJOSvzIfc4j+CBd3WN7q1Q8OjLUGshJEQS1RiqlBhw/aUfBygQXtaGYua
NOiIciTRU+5rR4K1EEPpskQIM0jjBLqg2uICFT4Wn7H1U1GwtBTwpkvqjDkfqZ/z
hgQavemYnjCuudPrQVlvgZIAJJGwh+VM/pWTSoTix7c1IYxw6CoM16BmzlyGugHx
v2QJ4sHORUFmTPTbDAsqgAwuNB4WGbrsZox/JSPSJrepirzQieF8C3b8lX9g5q+n
PkdrrtUxwxGdv6r45O385uq4EZA5K7UlCQmI4OuoM7PfwQJSnERJaUkjbF0AICBy
5YOGN4E9EuG2aHyizmqp22wJLBFRyOZvQrNzlxHa+EGXfsP/Rg2b1HPzvRL2ciKD
tCWJeO1QzSQqypN94nXw+OSIywfp/tTLYU0B33THOKCXrc4YoLJ1Vz/UD+iYoBTl
lTIPBgDm9XAp2fyHNMt1UTrytJsckDKPV7rL4wItp/qF4IZLDlEZ211WzeoU4bvc
G0jA4jpP6oYg1mtybzmA+degfOhFTfl5iFEXqt+vUNFsVPwoT4LFyY8zB0Tqes41
7a8/eoOrx0apWNu/moWV+HTJ5AjTSpRIfbboEWxfE4S5nrKRmql+rYZiwcx9AisV
lB0vP4zEUIZ2J+cfs+Ph49J+KE8yhCn8FA1ZzCVHYUTaZUzmbkCJP6eoA6OG3jHU
wUx8VL6XQ5ljDf220FMFRA5g+ovowFmzlG33HWRGGEcp2S7lMo9NOO6qHyE8cgu1
po/S2UTpgdImnLFjZSkttO4tjUj7xZOJEUEJlc2988yc6/ZkNoCKiPca3UnffrkR
hu0EDg0TzKJdtFSGl5MdwS1heBZjUwoXQhsclCiMOjlszle2UYA0pzx9RjzQrDbg
oxIItkR9f/3H12RHd3K+PcJM7YUWpeigTSJ+thKWfR4C4qGfiM7mwq2F/fYNfyU3
stGPENZbA/3AXKXDBOOpmGHrqjDaQdseAasdSLionbu4qsSlaLnulJAF4LUIW1Hz
w3iRS3gvNLOMUZtuyQ6f2FI+mgSRvIOISh1xWxLmyQ41Z5GzIlXDHS1byg4QLaWE
o+qwlNpB99zqvnK2TzXkvdWjIF6eJ+Ws10TrClxl3bXt6oWf4SEfyiLlgNE1jiIA
Ui0J2ZgVOAHBp5t3ClpP9EzZbvt1zGId07nzp3ajHtBiK6XQ0OklXo9MqLfEkh57
QqfdAzXiw5aA0x9HqPi7Zi6/UBEdIn4douh97XHPRfmDTzjFAWtEmoYYJB99PFl1
984VbOz6q+elTmqICkQTdvBPb3HroEw1S7DW9gH9HI3r/Y6H1tXuIrwORSvJUThQ
mv/cy71AULeA8Z5vOb1HdPEHW52RbH4iP9lEGfliFk2/fxVFtXFouymzdW04cUzd
L1dfIoBfk0TqAwS1/jMMok88pGlRAd5RbF1nQfKYrDdnIJ9Qvw60EDxN09khime1
jj2+lsJMnqv6nuUMlD9UYxSrm6pS4wIPPsKQdXlp7qW6QY+ncstKXPeQSIjCSxkf
a0YiBvmPZBPE2x/a3k5Z/dnTPh9szXVRSg3MU0jOvxRqhbEbg6m8JsMwiDbzKu3p
jKWlo6zrhp7MaJ5N2UbErAfXeNwUeWLbbwbJ3eIURl/LAXqh39WfUZtoVH+nesWD
rlK3Z/vbpnpXw1o++6wznmXsai7ERwklD86GF+VnN8/Fe16W3Klv46FnmotWGBdh
Gu5Yjf31x5rF9+8qF87We2eBaWxM1k4PcfW4whsumewdoM+lMackZBMnmZZ86Bw4
Fx9y7WuDuQu0++Sp6cBveCXMW/VLM5FabyFO5k0rPYqvMDW0P1DG4br/6pu1Iiaa
HGGTiR+yOjY7sYyuPqpRIqHYFI4RfZ3JXXfo5GppCIu1Wg700u/Po5lcJjdPlzLf
OcsjyFIL4a1sEukTrPQitHWBVzwB7zo9hYtJhU1VnX/785KrT5a4VS8a/NmL8yGQ
t+Yj2pfsvuCZO2P2JZ2SQYYJG3vNwEYdyYJxBtOwqjeqbkfiGxAmBKTS6NlNqzEO
YjpgAKrgnC7W6KY7EHCbqetWuNkbj4LlGhY8zcHJaYVNwBqKz07ACEjQX+0p88+e
oFi4m2Ac6M0+dpAMdL/MpHDtUfNrBPC44AzP3FzbQs66OfhTeJ3rHhonEua9eVQh
1ZxPuEoHGcAGp0PZT364RmjuAJETK4zNmDeyQeTQtMLbiJ+nnGt4sPRYWDFAn5yA
4ZPfmbKNJHV7NiP4/QCCeDUfBabYrdvxfLHXFI5gi1df3k5pc9+vN9BuBLQqbkXk
XspOn9rJH0ARDixaNTQ37i+t0nHRHbFpxBAcEH+IBvhfKHUXU1hfY7N7Pd35hRB1
EycQ+Gj9n2jXkhU8r5N6nV80eT+ae6huu2XUaIX088CWtnua2Qbbpf8caMFN0k1J
y0Ojhun4f4yKmjjiIm9+du2GcgEd98Rx5B/6PRHUhSb0HRj4KeFIzZDmvzfxfYE6
3ApkI8be2Zq/zQcRTsRiaeWM2QxLQWQFXvt6mzCrpy4HDLYu05kmOwRfI5ARYAe0
26RKqmM/Iru/fd/NhdFiLohJekTycY2iH1yWNtoEwo2oqFud0KUptF7/Hy4WVlfe
ecYSPQKd2OdIwlC5uIU6XKxRhTmoyH5Ezslkfrc/OBLJE3WSAZG4aWhv8ljsupVH
KgxPgbgNNT4zpim1NcaEXLeZko2kHgppFT5iZqwamqQctEaJoUHO/LguA28A/ydk
d9X3Sj6A6Rs0PScDjz5SmtOJ9mNbI1CaYm+XACR9HoK7b08qAUqaPwzBAHSLRHjX
7OykfF70I0zWFGNeE7y1LUokujmTi44qlkf9Fv8KMCUMn5hz2aXHqpKOkwUc32H6
oDwa0j6AaJdoxJwBUz480yXr16HBSP2LvIeFU4uK/YV4Z4xppE2vetRbr+uT/JRm
UQ04VqojgNvlcQ/UhlA1yqaOhjr+QN8rsYzcphaD2QUh2NZ/eoohMb+Gu7pXj5Wa
Ou5MplHr0L4h5IGNcw9C85FBt5MiP5Ez6iXCqNNaLF0gR2L0ZvLXIF6fz1QB1hRW
fsDwFtJPOlRfT591htSgsbfT7JbWxKFal3RUDfrhoDrJbIXm52WB8scETLM8cQSG
dPp/j6KNuuc8S+62kvMguI0H7tovxgzNyDM9wRIcz5C0GaNT2AZCP0bI3olApm6q
4uVFLxy9aPcIciFpjwMygc5Z4Jxc2Jmz+nMrCx+J6ZGscC1B+B5NRaw9o1G1staU
+eUPsSnXZjyfktBJ0zpJ7c9peSzU6FsV1zFfSkaURHTyx9QzAkugzZK5y7HFn42h
mZtG9xH4KT01ejf/AFUUHA/vOE0jsB17+LH2oZqWd7wo6h9n2TlKp7WKYhLyNB5E
gAJuUWLFyCaJxybzl7/8Z07kjSnGH1/ofkZSOF8kgDaLL+cgSyB3LLyL18K4RQpq
F2kO4WS19aWMCDX3tmDYlDNRrcsDOZtboVDXoi1tgNTgtf0fNHNFbHxqdZ+Do64D
6ckYGYUX1bdH8lyz3ZWvXWyMfOJHcj+tdfQm6Lm7MKK43P0Q+WgpxU0zzrO6ytMA
5mbnAQ3jrOoo/9OjDjnjBZjTEltyt+eg/mc7BbmGBDaAgAtOzACMesXayxrbyRlb
rgjR2IybCUyHSPLdJP6ItBNJYI9y647U/ih2Hunqao8Pj4FsPP6ZaGJT410N4t3T
YuC856QYlP6+skD5tClVdrg+IHuQb6f7Dfq4YEoyhLfODsoCwv7vTRzJilLEYCzG
8Crg7UB6pOmEswmi2WOiRe8GzsOVvACZ3G97teEEwnsaBgmOjeSvdD3+KWwKv6X9
p/RvVZ0lLeehoSGzv7afWiojAmIngo4q/GfYXubEt6QO8phyubmjum+iP+Y897ZP
v7ncenPKoayKROuog280SVLk4OT9y+cLN8tOrztDOOoN5OFO0KM4L4RXGOoOlGJy
FQ95VIGkb44i67rQWJZqWocbnOvPGJUXZJlOYVbXMzGpUJSEnZylbSDFlk0oJSo2
YcBxlPXXBwXtCUumiHRqRVymWUwgA3NlNdS0o+NXzq8fO0AqQoZWusG529fzxELw
QOi9/Yvsh6dT5UfgcU+PCOWaLSzySB40Fm1BLThwpbmY4a5DApa4V+uNBHaV6rt7
gsM9ajV/ypqp0VecVhThLHQoe9TUhtIhhTPjcBLpWWrclSIwDAhxv6weTCkY3lFT
8KT97O7Wy3M2M2biRNmjUmimnuh4IhSUwJOvoGzqL3PHk5qDHILe2VXUNqctBlp2
Ge0xE8fT1NhNQk/gkWA6XRVTo+JUuO1t32DdnXzOsaGq4aqefX2kVWpMKUGjE/Hb
1cg0V1E3V/YIDBxjWkI8ydKYX3Bm6Ecn0os3RA4AQSYd1mYY4xWcSuJVKxWjOgcQ
2M6JU5vQAdQqxof57wVE3nv2nInUDs/9pThjdjWub7AVOj1r1/6qbdPSM7QGbRIm
yi3D55p0gIQq8wv477c73he1hESAMvWBrAVPR0oUY80vdPomGKMQxSX9+n4Uc7To
R1/iw+S4UbY3WZVjevJvxaPc2oy82bXoLgjfRvkHrZoeUNiqBtbV7OzD/BA2hGqx
vjxW0JTh9EdkIKqzq3YHI0Zt71IF3tqWeY+55YpoFHxZjR1Bvh+RD2AmOlbMlWyO
8mIXMwW67QGbUFT5GJrsxuLbU+MHo38KKqpAcP8JA3CopxK/bRdNGvqsCz58StX8
8OWE67/AFoIQqSSZEb/mXaENtD7Ek5tHy9MrOj3qn1EtET5vJCbnzlunPrIiWaaU
gv3hLbRj7hLhQijahz44Zz/WXFUujDNvVirS8qGKNcg8p9NVfbvfpn2EFJyf3ZK9
A+yl2aPJpcBhO1RZnaVUmwJecYx7WrMHLiBvnFYD4sU3kdl02m1KdA2qo0UB0Kr0
fLN0NC3O3kESkLFqqMLAYwJ46eGDbXAQGC5aHF4IeEce2tE5ZaRh5oROtlPChDmB
IkCZut1gDqCUGrPRxbY+KXdpA5LNAqY7OTPXtfNIkrnazmtnNQB/OpVq7+q7Q+L/
OjTMxslPepIRF116u3GLi4Q+jmclsg8RqSOtH+H7pA7/HXlGX0xLqWAaRttcL2gX
kx0VUk4PbCCOVmUeTXOAUuzJdXlB6A0HqAOhHsKof28mJlD9TGlzodxKQQuFoTfc
V1CP7jw4wqf8ImwzmWgl32C5fSeuakGDPPz6QKJ/WTXhzaYnm28/fpEPjoI8mVI9
Y/YJ2muATNIWX56UmsxG59Dvc36suU7OFaVv+0ChRJked04LMhy5soSh401yHKy2
oBD2BlJ3Bl4iQ2k1ZXvJ8IMbuW+fA/CBtIp6MNKs/h3OSjX5OLUGS48gtuWWI1eL
cabf3N2eXKBtWsUpGDqgSWU1nh+s7V1oFhmoTXlOkTVOqamZD3cBpRSVdxyq6Uf7
ICWxabKF4FdL5RpFlAzfCU6OjDwI/1+knsgGxl/Nl1RHEuxOnJsEleH/fVubXqzo
CoJD27Yd1wQLQ5VDNG7vL16vbX1DInFS8/agJ33KyP9HI33C9f8ky+vcOa7qiN16
CpGMuj9FxH5NCRSL+uHh9Ls6bc7+O0COSJfLsU1USFf1u+tOUGeSyMrfeecFb0fJ
yWlmZqpztB4XP1ckx8598o52hL09MrRUZnq5HK1U6Rp6nLJzRv/0uhxsMrSsSSRD
uQJ8ixPpFQwEhljHoGQzubUgAbk3bUHcgr9yRt5Iu/o1n2wxUVj+ji4aO5i7oSzG
XgbWUyfen0lxss3BjiumbnEKno8aXHz9ASJeLwRwWR+N7DOjp8ciHGETvNwxODjC
RDalacBdSZ2XRkz6vFQjWlPd6WctjAmv5a6NTD26mI3s6nMLW6N7xLuUUYpXrEBe
of6Igc26sITvrlgxClk8tC/iVo4TCk6/JxnHwm57EZUnCUb92rdDWDZ3yMpWSwvc
su9vM8dIVRBqo7EbcilsfW6R6UlLukVa5bTxjQDgdAIw5CnkkevxX17+UVG7fyOJ
3ehkVrtvB798JJ1/Ozt9yMqclAmSoD6VvrvXWO//Uuksr1NaEk3LLTqULw2pztni
/R+fp0SWtU0tlKe2bR5uKC1JeykDP6Y8oiaQoIJBN6UqBevYGSAN7EynH9stugvO
Pc/V2xZwoe0COHKgwk3g8S/su47X2+W1EC1yUeD0tYigVIttJk1PrdQkt5f92i9s
BgNr92HpupTh7MoSpd52tumVFJjk7jIQxxyBKR5ajw0T4Mwj/aYE7BWeoInouBWC
y8QT1NK5EurnfBDCgu3Oo/9htupExPoPwi5xHIMXyG3QtGvSTLxEy+Cc1byeMXZm
58XBl82YfDYwZsKUwD8Mi6YcGY435Iab0zCGP4Ru4Vfej0rYX5U5rtfY146H+PFk
O8lHEAp0uaiWqzqoqba5arwvZrnEzKqg+ERChkGmeGF15qck+L0uHV8zFwjRszDD
Sloccp/MOpvWUn3ypwkixum2SchJXTLSgkjfRcq+HR7G4wCbVXCm0xfPPRvVU/4i
ipgTiRqQHz2iyRhmY8Qe5XqQAyTxgBqJAIxKmGd8Y4/kuOn09cYN+98rmtGfPFtm
9YJsRy5A118m5NPBF1G1Ln4ACsXircc8gO8Qbqhgd8oO/PhcYRywMrQth1QZhsNO
tE4MuO3YRDC2WQLfy/KvkYO9992nARRLPN3uQMpwFZayDlAoLNUtRBc38ubMG9FU
TE4Vp/PyXEaHoe1E49h5BhEJdSKUaplwjBlYo9fzVwbIBN+pqbNnJCb4aFQiu2vR
SOCXC8iRNmpqmPekQU6ANrVfsImzY9x7eQ0TajhtHcJXkEDBxMjLQVLgw3B/y6Ci
TdpOoJItu8QR9RWwHU760wOlOkZSSU7i46p0y07M4SPgpJf2JDttaYZAZHLgVQkk
RPPN2TAHs/WoKI0Lh8c7KUwRBFUe5ZXRj9X4tmbx/Kd8A1X957obmDix9vo79Uww
mSgOcEV52id9OKvyzuZNg65mKmRfdwWoDDhg0E7CeQkloEA5Js8l5OXmcaVzhJp9
A9g/S5cvo+9jakaNMPDLzZYypwp96G4Yee7V5y1FJE7ydtXtWK6H1Iyc2BDqkH3d
xULtgdJTKTRkkjK72pYo0ILhraJOqhMLSlPx+GnO7DpukQzKT36sVU9XpcPFqfQN
2Rqu+HElhlioR2KHSFbho/ajew3cVeOsDZyTieVbU/an6TOQ7qKQLNzW7tCdyog4
7w1j6t7ubLGKBl79ev+5hv1djTGlCieBRVHUEeVj1gE3yo7Ho+CA1k4GOc+Kri+I
A/0Lx4fWv126Y1ngnUim9hIt2lbSpCxNVV2fTvyAfSBLSHFZwGzgjj+pcuVTbyI3
050YCWlfhmcNHRP4XmL175J2eGE0VT3nOxT+Ve6DMyVaZHbs++eYIG28wuqbk/+H
TOiEsSCcenGZWBD6n+2v9vgSBlKeW0Yz/9LxVSFxbakD8+oFW6gD1J38L+G/NhGP
2YJ7eTYMx2Ih85m/gdoBgM/H0LirK8d+Ff25POjBj+xEThaIEGphwQr9AiIwnlKX
pM+yWW1ElhigMPazdYj/Z4fyKQzg6/fki/nIK10YvXCVRW8CfPZ0ZXe5K+DTtKQc
KqrIS1Sh2M6Zs3W/MGciiH17os70XbQ5oZbu/5GwQij/CazeNOvu1eqjVhY+YtlL
7CF8qRyOrHlyYV7lDd2OPDYbGxFWnjR97MEB0TV/+DEvuL4MXIiDawI+lZxsApdD
wPgfwnS/V+gLzsTJjBp/VyNestrxyjUlESE4uRN/Ar5AlxeXbUTUNMPcJSZXo1Wg
3HdkTrbvIx95MseNZ4majb49XnD7UnpaAnujUzA0CjRI00eceYGv3wkLDj5Lt2t7
qK2kSf4bIIv2stEeW6qcTsZ0xzt+dHSdQmtiHEM15fHHv8urm+x6/IiCX1ZzWmEz
2ILH4QCRqFQg/btEr96Ng2Nzotol/ZsM3d/YK6ocjjuFBupEomk8jlK8oUx72Oq6
tiiXHOMB1i0dp5/x4BMl384GX8owqTDMmcJ/sQvda/C4ivOlELy3klIRmMpzVBau
B7u8IbsBOJQyq4FoiI6sMSPlff84bj4AtkAVGjIh+lK2SKUHgs3964t1fgvpmAFp
z7IqeSTlaUc10HrVVYryWtugAY6B9Yh8f2awfKfT/2Sq6D7RtdsTdGLGPwF+cRFJ
UGrBm1EDpcjFwfDk+yGjnKzGajNh9csyClKShS0KR0BWBiPRImUnfePz6sVS/8Ro
rpRQBDlzfh4IvDM8oJzlMsG/FcqdbckYuYzNow8UbiNgKkM2SS28+1pKLaj1mQAr
MHtUIkRQpFfq3Vq/bUSUpOjAjhAzGLpreNMq9P+biE6SrNA1uZAtaTuwXHN0QJji
UjRNOSggkR/wQC9JB1C8TFb3Kbnhq6gKCEGCCXVYkNPnYmL4aXmiBlbDSgMRJSZy
ZBvZS1DtfGuU96Ns/1HEYedSi7tsttv7my2vzMuuGSG28ZhoPiLcGoxcf1TF9pCq
Z+LeOU4WUKshdi/cWy4i7cSBrHzdpGY7JAP9C6ufKDJzga7IVEiInxEDwI0G/vcp
9Wx9P0wEAUgDIujSDPA6H2zPFD7XukYaINHOFxAmntcbhLcO0F8Yfyzsa5ElHvIc
rMNLIdmXlUOsGl3DWRg7wVVFItXAo6C3PSgiYOj77CRk9twzfT2qyj8NtTcUtPL1
j8IqYz8KWG7Xzg1FIT9gTd+ga0bS7zh7gZZcAFY4NSSjGWolX1c6AcxBUAoNSsLN
wgRP/aNAQXUTKz3zWXRrNW9inAjMQGIDERlLEIlshXAyH+NKLw7IHarbiQ9uYdpz
Uk+D4+Gax0ibBLHGP58TvmuIHnI1+pDQR4sOayo3ZjLyLgK/0kxVhQUljbp3AISf
pO2ZSUzYcaTuOm3/DrkTyyVdt20YwAoTt+BvDqbHixGxFQjH3yEUmpohAiSxWYOl
E159p+Bp/7NMEnWXgh6LUYCefrnFrjBPsJkWZIZO2GMNS52d/Bq9roG4V2crXAmk
YKMH/rysQCwRMnSMawOnhPjrThtzKS59C3DK5OoIqFWFDImFGMt+To2rnyi5pF4Q
27q+Gah3JcQOrgUxGCutp+UPLiT0NTiZgVJkDth3Y9hGDEGAr8eeLGmyJOEBPkLV
mswe9eKSVvP9eAN6KRDJBHjN+yzMesJT7Jx5+HmahkaQGuRW+WjZYmUlJlumnWAh
3akJyzXE5DxlxCCZho9v5YfMW7+NUE/CDGjxb5zvRbT7pgLupZFmrpyL0JVxtShn
3wkjoddbmcB9xy7/Vj4QbktmTl3hL0hNejS3RRrYkVQNBEjUcZutN9xQKoLJ5ugu
dEPKjzPRPFqLoeDTuGUubhs4WmgqBww1GhUKn1q+cf2eKKNaeoXDNh9PKSZJA7wF
4s5OS4K1vD23viaSf08dq6+rZmIF+Q2ucz8k0VLUpuCEtWiekXA6hsF9kROtFakF
wS6J2VgqKc8jbhpRhWDYELOvHtUS1SCbehce68C+fGNCFAPkazRUK2sY+3e7Cyvl
HW3gHP3jeO4B8l1R/c2xJeOIpsjaD3VzX0IlDAUkjUKa+P+0tHhKpdnT7aZA/lrl
xOhx8a34LQo6w3OGjcfkwKmOCnfOdfQSXlux1gbgcXHQGiRGFZWh8Ft/065oSuaO
UUYxJqQiUKU4Csq+sMrY5hpN1rIx6ucdimCwhq8wfW7ABJtwVx1aILcINuKU7e7l
ZQxAmb+RgttrOMRQQoLJW1u4J2vrZVibSqpYlGADtAk04+2gUxmCQxlRfSMa5UOR
Da97P/SsMifYgk8qF7G9rzsjohPpmLjhGkeYT8flEyeipEK23Bp3n6pwzOGvySBM
XWiUSXqJxGQ7hxxg88WmOYrEgffFEQc+ayn0EoPlXJzLiV4Ht6VCzWJjWRNIEcaC
d1VVlWpP5r7rg/iu1W4VPzuifnVz/TSOiefe7tjtTR+i3ta+FH8vJX6JZushOyg8
0h/aXp+M+9lrE3S6iVA6lZw61LOwbaalCAcCZk0hwf2ytf5Xmdluqo/TXndwnsXU
IHPHdyyS51qcpb5+SxviKvN1la5TUJYTvGzPBQB+CaXVFN0TB15AcXREIVlhlr6B
eO2ngsS2FoYm/efIOYcPezVYQlPw0ORSIExCaKo/GD5Bm6XGzrmUTQNv/xuIC+J5
mZB242ge5L56ilOrEOzSvDS1jkqJhuG37uebIBmTFAFLu9MDBJB+Zc4llAbubFz5
FKcegwhaW7KsLd758rZOIChBDIw+O3omJ6pB1XQvz/SzMFoKo0mgDU1lWiUyIQnV
gHJDLL2dDgmwh5cAtCzyVv2/bNIEkYK/aSJZh+jO4zvhnaB0wAeEGNnzZ0qrs3X7
M3q6ujFmgPRi6K5HJtR3mTVAkFUBJj/5EbqIGIzQgDTLtks41OKNL7WhbC4AS7Q7
ALAshElIcs8dmtPAGX/YwSxEu/8vkH+BejxBrJL9BY7AFwSKPCrYWvmixkAbBi7n
04L6hKDQ/ZliCrV1TwF8XDdkXNv782//GO34uZ/ahKuZgs0aPcrK4WJYCI8W7bEV
bRcZ2pN+h0G4f4+8nF+Va42vI201YB/L9dza+DBBtrF0orNdcAVx36yARH2zBhD0
EwYLlPSrvxYtkc/IVevdf5ZOpmyIcw4LAUnCPtb3OIhBjz3kJNXS+ZYq0pXeAJSo
YNgN6cdnEMA7nDtsH0mFlxnTZAsH1oBlRcgKzgH+hsVxKv/lhN+qMpwQoEQm3zpX
LqsVzkHpcua66ggXXnkssinQCgQQBeODav+thgaa8okyay5mkHjmXMSdAgHU283e
4OODsq+aARn3igw1ffaDBjC2EEuWFENr8D5yRWHQoNYWReCq8kduIdpKW+aHG3nD
O+GdDHTEEgwtvZzX1cll0phVyY3phENVyI8cfwE25/2CY4yxggrCPGdxkrKVDe0k
IoaUUODPsWOLrY6Up2NzKA3obMitM3FfmUH6ygmgOWJ1VziGfvEKOgbSmxj3WBbZ
vJ/Wy3thROIlUL2zgzWhunhoOrrHLiBhIVa2F2JBxzzrwzmY1rNEeWCJ1VnDBOJD
U3KIRBQ+0VSDop7bhdpQfDvie2UvnbaEYdWRlgeCRXRE00n6qWH8GyGVh2NVQleD
+x1N8YWyqDi+sEWWZQ1Jv6zUdvohvVzmBxR83f9T0Lt+92BVlaIIWLucqVdBovnN
9Mhi1SVkKjkgdr737p9WKaLZFlIe8IGDNu+5jjyhk5eBL5s3EFzVNiH6qtT44Y1q
s1ZEuiTk8AbMuBdM4Puwb6szIgJHTcDhdVProyB/aehdSWpoNDMxyoCjd70tVU2s
4zUDwaesEkUmIJbrCWYqokF0cjqem7Ck//FoQCilNxHguIiAN/8AOGDoDOP3b/z5
eMUNWYweI953qW0AtIA1W9fLZAjvonYQJnqnq7zRCg+sa3wO7syuU+a5uDlCkjDs
jlcuHOT4nqahbsjLAwko+6CnRqlRxIcDBOjPDyXaNiWOdTC1XE3Wt76UJQ0HaATL
1FpDrpEWBbg30xt/Qp+gTLaOUAoooZN5TTBP85zSP4jFp/IePPOdT6ud2NtxY2Lf
ULM8oQ6WCiAYxGujusVIli78enGpKkRCKyL9rkTTtqKz/4k3aSwJbyfR+4lchamX
KhN+R1nXhhxHjCHVDs42B9hJNhGLvb6sbDoHG4FCUV9rNtD0ny54zj8p2gjtESKn
kRHHrR74QZQvShQi2TDUiCz/2aDOlDs8Gmr87YXj8Xe8JLYLgizYccixwii+YKte
UrktW4cw2gzAYeHo9kokzzrkvbipPoKL1VjbypTpzsDBXhmV4J/9/rbnfSQ+FI/5
UfYyhffcqJcPEw3oRC29wsar5tsJEdEV7gKtAJXVJydexm25TQ9zm2lNrp+UhK7U
sJar5MUcVqZbuPYzizmdEoAo0jBmxw4tMWX73bnImQQ3e7seQrXdE7iNBoltdgHy
qCB6GN/XUAfBEO58fv6LumfH6Ftwiq13aHgy+B4QpU38aJYs/a/1Zm8FzHtaqQeh
OyJingD1v1W+3PXYGkNeiYrZ7Y1xUveSUU6g1nXd8lQ=
`pragma protect end_protected
