// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0.1
// ALTERA_TIMESTAMP:Thu Jun  4 11:11:14 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c3ajPbBy0XemrqEz8e/wDyjBWbk70quUyZtn5pA74uxn+tBxe6L2G8IvBDDjPyFs
GjxwQ/KWBBMn0d7aCrR4v2qrHadMrXdXDzc+TaUnS5CuNr2XkTclBWKSEp8zleNF
fEorjlAfHNNqaAOs8uCx2vPNdqdFoeSruJjnRq/UYPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
LnEs88kN7zDNrxPm9CiawB46D4NSuVbIlvNTRzWZvMDY/8io1E/Kowg0giOpMohS
I+EYDfqWYLTuyfOA5QkCvwWXm8P/QTPvd/xvHpkgbhVMKXte6QWlBMQ1fqPDzfJH
r+EISXsBctLKdjGzfDkfMK+sAzhuepnLjDYlJ+Xury1UzUM4jhGFRgUK7lW7q/7V
ZDsajFzJjTXyYk0hm0F9KVXoU/Rv1Ts6rcXEPEA0ef8ipQXuMxuJsXPhBVQ8e25C
DaoqFo7PSlhJcg+XCVKykOSnNp+F3W53pLYf2v7mYn+N1bNGk6INpzUq9e7S+3aQ
yBp6FqyMmm/Umx4jUDknlRVHzH9eaAu+F7ZpLuZryKeN7WydWaKUh8eOBShYkOSv
GYsYJZ+9cfkDou9j23xAGUteq/sBXvN8qOEy4Aj07BtdhJYBBMNtZvndYDmM+982
aW/TJ3u9aEVAfZjJsUGgqCmrCpRxLPSKxD+ApjcIhxg/EbKSYItIjm3SJ1ONZh9w
0xjqhII91LjbAYWLVza/wBss+Y3bGAf1JXAwP2P6uOOfUutbJoooKmnsJfM3vCum
f10UgvdO8X0uOYLGvXeEXk69duTbWk6P5NkASQ4wdqb/kYbAc9xv4eSkE5ReMi+6
xGsVznp/bHln8wiFjjZy3tZjGn6tg6ND5RJmb2XdxdzmiIgx0ZBWATwIGPCrLFq1
nRnB9mdqtJ2pd9iI2icVNYh6vDIC0LpgZTFtt0aEtgIMWmP/T2FF0nE3Wfpw9d3K
66r0101PP+HoNDqq1rPI/vMepLnL/y4qR+WUSYr1MAu4+DH/5CDfdMr7o9XUycCf
hwJJ8n0XRxkRG1nmlZ+1qrrKR8qJCXvIG3KWXVxX/b50nIg77uDlH8AXUTx+G9bP
hG/Q0WhpYpO5/Hls+tAbezgKIydaSggFIZcO2+IuqWrrMu2Z0zmDg5pmG11i4B8w
iUm47rDUZ27ksnFBrf7MUqJEn88CUE/0hYgO3n4altQ8fu6BitbGRXjKkG5YGHue
V0MCl2KcaXNm80LalfzZtTiTOXplh/ByYDvkLN9pm6h5zj0SWDC1M+peRyhQs2wl
G9FlAvoaX/EIM7+MNPV9GdHLLiGzljxQsGhLrNx5sueaXU0091CfeLS/l3HcFEUQ
hjFhp7x/lkLnPa8LHaikagzLFJBgEXR6eHh5j53FQ02bq0OTNrK3NoN88OqZ76UA
dLnJ6qbvjCAh/w6foqYJn7SsegWmVwVx6nVsf1ecbo/Wd6InVaexPEqlNgdq8Fzt
SskNXUJ80AOGPeu8eiKCrcmNbjXZ9XKZd9DbWp7K3ReMpHiAgcTgGr7t0S5S3fTa
4YT7VNiVS/0IBB3swn/xMiGF0827qZ7zr2aebNB7cVaXAck8oPGC1aVQOYrGEXcz
DKyynGmanx0fRb/CjFqZ9uBhEYUa0sK5nhCQL7wTvMddoSmY2ej2OQe2zEStgH2j
gBc0cAxHrLDw2n2H6A+hh17Rkdl1WnIq5NYCMWEOrl8/T54j6Ugd5YbcXHmlmkCs
2fTQU4xhA0SC+UMDuDbHEhBD8shcCG4AM7tla3wAezl52Q7TjILl3JN2A1X4O8OE
1bZ6eNCouFYf4DS+VYj21MQZic7OxGJ4tW++0eHXQIyiHtT9dCNSX0IRr4v9H/Hc
bP/qdQDyspdOYcMzg0NsTKYbkYGr7eqoQFY36Z/4iZBjP5Fw/sk9taaNfAc1zMar
S8bALJc6wafAfhLJxY948BpwMzRG8lVr2s1D69PHi7TAjf0ZMt8ANORU/AByYr/z
kEWnHx5lepM5tygzZRsAlPqSjBM/djnKFNDhrRE64GQdRSt6KYH/WW0ldJFQHL1+
OXV+P70QBbofBChSKU+nzvBhon/NF2ztDvmCdisZjNx1a2tWI6nYKElo8ElrXRQ6
BOKnvFTTRgpQMxHUxFbefizUxLktqEkZmEQOOL4/+GIG+iHl91Jg/4RKNH6O4DUH
/dv9UWOLrpLQ5EODidrYEI2ZQskiwEq8MHNKs12uEZMpHhNWBCZzpKGTBagl7lUj
SytlVY9fvnuJ5wovGtPtbfnEEwQ9shYfUGdNbGtozKu369iWk0Kcg+tEEdME/KL5
jWM7iotZ/DUsREmbP2clPbMFCZDSlYaKqkT/loaxuVtiuek0JqlIAcNWIc5TZQEd
41hEL9AynacdatwW02wLXtoEHrAmDPCRpyTs7anFc52RE4xPUCPoxxy/GwpOMJSg
JjWxHQZ0p275TysCFNdSNwrsi93OfFvWFoBONE1H/cqtbv0/baEh26rrKPZ3rmLO
rhPQyZeIZ+ffBMFDsfR9P5ZYOiEUhHHwyyXma/xyfSvPr9XfxRqFu/QBv9EQB6OT
U0O+WzHD57wdo4ca4K+ePebD1xoBQtRBcPLJVMqDYmE4sgAxyfPgzkRVBifrf7Go
rkmQlWyPtV+wicR3yu45zuY1Ziy/+7j6hi4eJC5teD2Up1jGuZFUxeCvBw0EhLDE
8u0lsW7hqqny3YA8SWPiDx2Dq+C05/MH0xq9x4ok8sgc6RCt5jp/PG+161CvbSJD
5TAokCd1VJ/7t68LEp2RjrpNJw4ao0dAur4hWTJ6ErJ7hmrg2KiXNQstjC9ysMOs
iBK5QcQ64CLoX560Z6imXvLxpL0Iwfyn0Bf1f7irbTA0rkoGQXJUytwKuoQl9k/C
LIfqDz6yIyUyWh/Y7pAhNXP3YcB/cTOaX/bnvX+FwkoFRjVuB7a6Y2QryTGlEUQ0
kFNyDo4hS31MvbR7wMyDbRe7vnzssOVMGhNd+Vai8Knxmskv+TASFBTynvye373c
wsmgHRovHUmHGu0s/VI/vKQrhUrEY6uibyXKJNUPuXrieFXj9KwJeYUV8vcQr9JD
4qOr5keonaUbYxS199CgZNqku7qRLAt05OGqQeMZnnT6Pi1Bzwii2uxgTKVZ4vYB
zITpUBjKkQWsL19ty6jUHig6yBKbtfWZ/f2x5mgDmy9CJuYTZjcqoXlEZArHJ+mR
DjtYuJO2Dwdu3SjwJv49LYP2Ky1Ite9fag0K6KGpHbdwK80RlO1WkhW+KNLPXbiF
F4t8uiZhY6sD4mVl89EW4+awaQ2AoFlwxE0pv7KweDk7gWtedVV5TA4jqtDi31bY
cwPkG1CsUks93VxF+ydSSpqrintZ+//5NvAfiK+HbqO7ROzdTzDRQ8FwuzSi1Dqp
j1xMHeXc4wMy1JPrMD0XAGObvXByHWjy1uFCRz25mZL84uRkyNrk/DYrZb0tVEkP
MFWhtMfySL8mPQRGKgRiVRQrTdjPHBcAD28EfVShRh2J9buOzhXlty0+AS7rpcWv
wU0QH3YGDxdv9LWoWJE7lgBKHt5rwda2xtdNYjJvl+BCqcwpyrko9m0E87iYkzVF
nv5AVWdMd1iG7n4cMDjZKUwsgPUGpHlWEYllLhASJMnny3meDqde+geo7wE8whuh
21it4ZVmk/cd6BJXZLdbGFcx/jj0r9UOZ8/HjOc5JW6DPo/cdAgvFgygo7wn4C3Y
2ptHEzLplrw8qg5LXjcK4rCUQAVE7kotcBzYRflTUfqRyCALGsjX0WW5ZZldy85R
VgBULZ7vSvrFXXzpCSA1R5W8LHW4MK9IrWNvA81GEXMZFE+0aMSdXQ7uq2vhLsPZ
YrL19tHRse3Mb+udC/ImKc5+FKul9t5SCQa0FEu6XUrhv1+ZoC66tx4nkfuU1ePu
I7/Vyp6RrxJGQfMB9Z1M+OBOwY2EDlYinPf/gXc3POdBUomFAFyf1PggVNuMQFAm
WhjUUPIBqx3R1U5MBYNaUUDXr28C6veeeltBIjiCm7aZ/856XJnUA0XOcO5GBcgt
nzYu5XKdo1ntW0sjTiPuLpOrlgaaKX1QNcI4xfuygMGSm8hyNWgH6hwRhHklGiPt
idxwKo+Ewv9EUXTCrhQ9v28OD73VnHiJ5QnFSINt6CpmmpSSN05qkjTBJ8JgFiyg
lnGoeqpqED5AEE7fapBFPZ68UhHKHdBMmQCR8ov22QH878f/qOtWZUyjB066uV3E
r6/rvUZVNafBbxTWTo1PeiGXT8Eja0c17iwmtyq2gQ99hXM7GCl6DTgJQxcknANW
K3dPg9TUyV5u2FRbvsSiymssyIM73Yn3xiV5CQCfMNoS4JX9o6F1gCK3g9fnnGuh
A8TCqyFxpoPspdhi7e3KwM3YxE2vMweB3Nx+ftt9J+2i0HrLHnDoaaNAxDhl7S2Y
vwMH2/pm7R8caR9Zn2NAq1AOBXNOHPIYWXZi+Eh784GfFAjqhATc14523xhMIBf1
LoJDN6DJW94lLRdRNuNjslqWVkp/7oXOc8C0h8UgMX/eBokeE01NYQaZ7vaRJtc+
KG2Qo454LU5bgnL+SgY3kLeLomGIJXOzXbV8V7snJ/hAyGDd3qSV3ogGUgi6O0IK
+Tezi1ovuBx6M7K6PwwaCYSNUy61L1rQy/ZNSiKGjyyQMIIDVeP/OJjlVsCBE42Q
bZbU8ctwK8TuKcWyb+dw+k6uP3O5mVIvD5UR5QQoxdLpxW4MXtKF30nv7eD5cBuw
6F0nc3VoQ3iSxlENB/Wr9GCOmyPT/aK+gGubQGSshe5ShYWHcd5yg4v+BgRNZshK
dxlOon/10xELyG0BU+ou8O2Bes7z7cQlLyfJRSRM9of3p9hVAkQ96B/5t6wzIncc
wQ5D+B5RnG5Wth2V8AMrVnpX72UyFSG9l+35Axq9g6I6gYXd0kJ2aC5KF3mIKFPN
UdE1E6cIffVZz8Ecr7WCmciUegwo3nj5arYMjLb4DpJ16u6o/dzoHH0X1VseGC4r
R8D6PvjmcDkxmAlvzmePbJtfHtbaK6ZiRNKHRaE1i9zx8+kD4/bOgFWqcC2pGjER
EIF8egfuvevw2B1K60Q+c3/Ujnixu4c6M5zvBqGSlWkEtQj2TFP/PwajI+e5WYQn
XrS3TM5HZlQCM0oW7zmXkPhckDnTE+5U6KxbhIfDU4IBet9lO4gyvj4P8JPGaOGm
zNWjQVqibZICQyMU+YiQfPGj6i76IAOMzp7iaV2pnDMmRRlc9ZNAn7dglp6BPWQL
8P8x0wuEa0QmY0R7KVOY/vvSzh0BgNMZNrt/vvBvTAy+JYHe6UGVLUh0gNdD+LxW
YNiEwWdKBitWIM1d5UJNO2Xh8bWrBUnWy/BDwsUi4fscnGbJ8OKjxXREDY1fU8kL
3L+9ZlprXSUuMIyV4wNbmHG560q9LeU0+XDFTj3+8OGc2xkJpdMfzuCSGkJkyjG6
59+V2A1JzB5BT/PrWTc9hglMKywqFx2pbGTNrwAs8rxDJ3WYcBrVn3WwTrWD4z3L
REG+IGX7OgZ4wsB0Ip6aZwijzyDXXsB300+sDypYQnYRsFl62lwNZIsUp+AEyJ79
eU9Lb5hU84UYgK0BvaPMwkLv0WJvZX57LeN6kuMBIanCElCDwHaT7lND5R2zTmZI
A+1aCRVVKTe0QIp9HFnsvoWOED/uPXpeXbLlizcwNHxxukmFLbpIHHo8MTp63tJL
3LeHK0kTT36t6CP9uOUQk4rcXjSUypKLwwRqdLkKRqaQ9987xtXlyxDBXaX8IMdT
OV9YSuf5MuwT4GdW9dVC3sdwGezXANvHDGjH3Rlq+2PJdZ8s8zilg/yIVUdPRVMd
stDZQwCAMDGSQFVtuwmtDDeOAnQW19pkp6QRp1yTIrhehZvrVZFlr9/PcqqXYF+z
pAdj6FAQUV/JkDava0xpZZ+BXOlkzMRPGMpDdH7lJ4q3Eij+KMUW6405PKB3+MFj
yJs1+NroDZPW6JPinbZv80ScClIcDc1gmnC8ZAkNe2yIKdWzSoH1pyJGje85MJkx
PBjhO0WsXJlexB3zUlAynFLrweMehqYyrI8r9na1nurW6XcKtF3gbN8jXnTCwSHS
7uG0CwhApPAiPkX5yeq7p/8nRFO20kUP9AGIW+D7zp027H+rHPjiGt5GLZssr1QC
ptoTnSzyYraPSn1Zkes0A/RrHi16ULvhDEe4jTQ5/ug5soIeeYzafxLE3VhNZ3Wh
U9qDohese9Q3RihG7Pf3++b4KIttGeuRsmzOJQCyiKjS11V/0+FoJ7y3qQ5ZqvvQ
66Ncek+xMdDr0BNpTo5LIWLqrRMtLi6bwJdfR7sTadZxyCQd5nY6YkspDWKYf4w3
z7ELGb+cMuqMd32miOKltJDrUqKvERw5iaLFqXVeDebU8QOYiqHc644l6rXt+Uxb
mC0vP7TVMAjpvSsJZ8z1fkXIRCwRZu2ygm72EWnj7RnXZju/HEurc0+V1EvStgys
R/c/ne0XlN2YPo1g2uNGDdnOruA9RRDyUzJaa1SNCnGAwqfclm4fhV6BOp1aDKv+
2wE4vq8jS9lFW5XYI9aFMkGHF+toov3EFCYNBIeS2u6xff3UF5seWPThqRjgOvdK
LBPQHC/kJ/NrI3rfezOQsnjGeSz3uJOck8ZZyLgfJDbu4q/f6JDm8Ym7jLky/ZK+
LyiPkccs75yZq6kDC7kFMhC7CyD5kATFThlFGRS8MYGyZMynuYDjQtmfkbDf4E+j
/CSR3fL3bxTtqJMdNbbdlG7oJiAGvVgveGAQnYEcDmbyRVQdCnAy1psYWWup+ZYD
LGCIMtTBB4q/1p0+S4GsN17EkAYMSYM7Xis+WN7iu8NqWfvET8kUvBfFG3bR3vcj
QfbeWHg7O3Sm4W6M261K3uHv1mHJA4V9G0Pchp2HRMoCfwcjUWaqVZLjF1qc9UiJ
Ecp4D2dH7hOYQ3Dd5apvsakKovWAUaXmiwheLeaWMhxn7T+HA3/jcrWXM5Jc1Z12
hoWXYvX2C6pCjPZXzpkcm7RqcgdV9lUCyMweewsgk2ElErKvT/0JFxJFaE4t7cIt
t+V2ZT1yMSfQmWZYcsi8PJ4BNl/R4aoFailQ3NAQCwbgtb862d3G3xcgxB55XlA7
f+pXp2fFN6Bk6Dn21ylXKeDyNV1FVMIAScwbXgfpBM38d8FOSmwiInwuuxiu83yf
nNmr6FFvd2IHvrXyF13MkCgC6kQ6x+eWTu7jBi6qxyG7qQTQ9mEvIaS4htFmX8ZE
L+jkAEvKR3AOTslrJysT+Vd0J5wwS72D9L0gnLPDZN56bZJl7ZgYhSJKi4iRSo1f
L7nri56W8FeD+pdN2wIIyoL9u89b757wfsy7AvIGfi49uqyuc7NrAt99IiRIYP0s
FBbzwvj6h1cEU5YKyzDi7iS+XyNVeQ/GqmUFXiJnKOMi5mM0QP703EX05iNGGOuc
f6WshDAd9iG1foED10J8wxrdvSCgAaXo6OyZ3AfRuGUD1UsbrKdrHNjA4rkb+jtP
PN8l/SUx8XJjJ/C2JNEoK+CFY7Lrl4ngiLnfi6KmjqfTeTzZPppcG6X5ZkQNpSYI
4iWgrJzofMWRPHmCq6r7M3cBWcilgUkml65n2c6rHKAk6LsHZc3HyvKGdBqbjGAo
UymsYNxcClEbRb/jRS5MBQbdsS3o78v4LkdJj9BcqgWsMs+VNToD1ER8TLsXEIJY
sY/lGrCcu3TwGWdtUYRUQiSrRM0j6ishtc5ROViGb2AVYvWSfaYfDa5KpT4dEyPD
DIOUdw8M+wmrGN3Ksn8b7lpWaX7+R/apKdRq36yImG6lf0oWvxXAjgJQHOoRemch
sFEBz8e0r7+ue57+vVjRevhimxPzdco9DLZW7xrppKW9sUzvyYD8kbrfoinekuPJ
5foSgBZsn3PVzXyAnWOI0GXDNK8GpUEKSFs6wBGBdtxIKih0TQzWcXFhD6LnlWJr
qPdGjHLJs68qrjPg201vNr3TEM6G1SXI5rnBTettjWe2DyszUfGQz3rntHOGcK2P
U3GGpu+u/0RqptBh9DzqEay4bGFIixPwXb8SI85tmnG4m/fjeMsT4t49g8v5uC2l
0oRJ2uizEc+yj7pPG7DWZsoaQ+k9FPt+lFPyrCNqqPpW56oosbtGPsiekpWhVwMc
v4+ZbEF+slUP966xpwyWXsTJO5X0ZRhc4VoG8gwX3lcOzmaYtT3BKI9Lng3bFi+o
vu/+tivinS0rc0UB9MiK8+xkWz8gIYy1Cxuwe4H1lmZ3qhbQdF0l/Ye84ySew3hS
qx2KAO+U/Tphn+uQXFxrI8bWzoOytuDUhrnW8YWQTuW1CeDALVtPO6Hr7mwvScu9
L+SrHZn43bQMr5i/W6ZUeSrkCJJJnocjZcZk7l5ug4/n2pTZxJ+j8A4+nrJQhzcJ
HLJIddCujnz8IoEFE61/iN/oIMZF54OhU5BdppR1C+hV7QtCVx3z/MaDuKfkJbKS
GuqAD63m3vz2zhpEp+b+f0jzVeuLb+MdnJsdGC6zCL0tXhuvO6fWEM/MnJbLB9lw
70eya67KqUfKg8Q97FcjqJNZ9R/fLrjE9HFs3kNHlRDLt1mYFJ5SEcl2leXbfrLX
20ARzqDjRYyG7L146xrS+N5ZlqH7ZwLrEkYnzt7oDDkKAWGKQDnzckeGzs9wRKrV
9o/dWJRXP/L4XWYjEsBP8Ceo5IaPfVvngxTlZVe6eK2oR29snttdDdzW+nTJ9NOG
JgStLCUWSmDTtN+BuVlDH3rtvAMDC6JbteWUeYIQ9IyJ9pD5tyHGvtbr9z0vsHOf
RuQ1izfSvzTVZC/uZwkyr1fgUHYdzLHFRhtuntKzYonu77v2Wrq3hztFQ0VJnUJN
a1GdiItrgXbD7bDjDIuYqHeCJohzyU/fApyN7Kvlo79uV+JtRvrStrRVyxeNjyIW
9huQ4dhy+aKSIO6lSu6yuDcq4ZejkopqkzSW+1Xa2unVLFUJTBxF3d/l+7RvCLVr
+sWzddZiQUFaN/3dRK0cfSxVtFei6jND+datpfCxSORHJPBFcSicZBT6KBiwtZjk
Dp9GUE50EaFHhpRWXgG3vj7j5g4DMbKLHFwo54sxlxblvNcpb9iwFji2KXAMM6zV
LF1maoByTVM7+bskARvMV4mdc+ozI8A0yOGUdwn/7d7938tkb586DZsMM2h2z81K
wf67WZGpyKjFfoCL2L5iNdob//jXdkSlXVR9nQl8gR6aB3MIETcHgdRdHcn9xMqd
+QvdH+exsXZJXAemCSiqFU94HcQL/M4TR/FQXpZDAapw1Io8yuCuADC8Tljhsld5
LnF67MCzkk4aLI+rGQHVdNJib26j8fN5tpAOA9IEh5Io4HEGBr9dGPJq50UFGawg
Z9PXub/GrgsTjwDykt+UMVQf9Ma3xfyKsd1JOd+/Uyb1VupEhU2c14deamwZJb2D
ruRZ37/DKsYhL3O0FWV19RJAGllahYrSssex1zrOsfeZ2rcWzK1+Ll2SEe104K/S
Vvk/Q0UQ2no4TyZoagtiABL+VkKU7D6unDY1toX8HHQq5sJ2suuqPmcYRNJUgtZk
tezHeetCLnmOC8pniVOiOsF/h8PYZIpGeAs3906eMDt6nuzbF3otf31SW+gMIyI6
lFDLeN5CXuE7Sq/QqmodKz7fGUL3RGQrz3HAR/0yIvmvKhbcVSSdtKKAVyQT08L5
7bx3j4SOp36rUBf3vZf/hihdT0WedPcWJ+KxqnyvkCAiw1ssoTIpQ5FVGaYeoktf
xCWg87gKaRFkOUL2Ib7CTxTnzpb++WaWrrhsb+nDTwCIyMoB77k0ZIMQa3bYKypf
cZeE+MA9ih+xwA/HxUUkOKf39XVD2ovl+AaM7zar3hVaXVECrY1tSRqxU4l4flWp
9S89qYI/OlVnv40/GK2hzf43RhPsEQeB+ia+Iin2arCVLiQ9VXswexJD5SGuYqp/
81CRaprQWiPsy/+0p5Shx0VRyG7Y/rQ6miAD24JrW9Sb1+p7W0cTNiG5U/LFmhY1
RxjANIrtBzmOl5lXVE1O1fhQ+KoduNxhi8VN4BsBw+2rYZeciY4MY7t+3PSW/gnj
AtgKJB4ld2Lkp+c5sB5a5zddBaWT43ZY5El3B/ZS24CKjeyeNIhFyUpBW126oMNd
zK+g+JuN6ldxor69p0tv1xauTqg9vgJuNqwlxx0RriisAOHOnGrrNpeHPXn3IMAo
oYt1qHCh8npTQvjP2ZqLZ0b7egLRJbTxvQWzBDkXwF41Dc7+E5WK0XLA1j4bDT8t
ucOCFvhzdALrxxcrGHyNaD1a6nV2RNWcwTWi13hJlsZZJJLg0LNDUDaJvYQ1BSj/
I/ZJ6YDXI2bWfuDtdJrWiVVv4EQqXn0uq/c981cD1EIVXCiKUwbsqUj/i3WNbFGz
fx7GYiU7Ss5uAY4/fPAJUZ4UvJMVW5LzbJ4gRn6QmaygNhVRUuuz1mxxAaPEMk/d
K8v1Q+rHrFTbvvYcp5jgVzgAczHp5eG8JfrAikVeooyJ2GaJemWhwoujiyvvqvfe
0YpnboD+c9ZHd/Hk49QNoaeunT9lwzur/x7Lf0hgB3Yp1Z9dv1qadJ/fKlrKetmO
tFbDGQKj9++BylcfN46vfAGbgsVAS21Rs/2PSxbWiaDR05EHBDzp5Md1gCZU6ITr
UBBjVePLtKR/whGkQD6gjMFQVfqtePRwXIENOnsVVFZemdvAsWS2BPOt8dZrgvzW
ulA19SY0/hPPCiYG2DLoxCVdFlDgdXncxP4A/tMiLUu6CW4SGN7s3Y7trXDjbBHV
zHAiy6YiH/QDcFUzaf27aG3m1i7bY5MOsOT2aPQoz/l/GOESIgKaDhoocDi/G1v1
Yt24UbufyfJg0P9WQtege7Ei9Muq7aqJfTEiYST7ShOyQ5G8r7RZbvFY9pxz1oS5
EeB65LIGxtV0xr1K5Ufe3DrmjCx2eIjtkHpZS8RY/IKbRxOrDWveYPd1ppatko7o
QU/dGv7ncdsqJS+zAFzBoz6tEuIdZ2fDXQVjypnR/tIdcBWrSZ8ulSe9PG/uAk8P
/lTYWH5bx+tajXFSzYtiP13pAuS0Nyc8s1jS+yKnbaY181jhY3DxiHEAt+Ru25i5
lrxw97T2fbgbjtJsIC4rEye2ZLEvdTNMSrm/7Xjsqzo5G6+1KyR4D07xKf1fU1zR
Mju4QQRLydw9l5BO66cEV1YX3f7Dc+hwd1cnFFsTrb3MCr27HDz+sFtEmgIoAoRD
TzevQbwM/1HJBiwx5CMeeGgKtZ4vchxlu9MrbhM8Rvx0nyrmmAxp6ivwUonFZBE3
S3sHt1PELEnwgucz0GcQaWU4ibVHHIf65Y+rUiJ0uFm6hllBRPS0Bg9GGIlcSFAt
KrsBW1CscV5iRDSnIy3WgdN4gxrUffekiLXKyX4vW0tW3C6UbOtY06QOQ42FZaPD
xkLxPWmeVsumCqGBR/zGykbAqVR7YEL83JIKtpWWYmE25pNDyK/xKloG+nvyp6Mi
PRw8Pp5wGngiRpXMVE2H3j/7NcxHC8DISRd2nl+VNDRdBR1I88mnViQxw5m/HlOT
DdN9pZYfXxuZeQMSVaqZDhcJaa/eWDksdqkRcz6ta+nGWne227stWf77CqldXQc9
Z1HbjRt+1c4PnxYdlEpLyYFpZ8dezFj04QhmqHElFp8j5buNXhtSwOUnJHBXDKKE
mFZZd7cLnSnqS1ZPtP/eAhfnHmU6cu4BpIUTsDFt9KYsKYf2UoAI2PnU2vGlCCfg
CJbv1i9wWvmuO5761vCDV8PjgOPsOzS13rLE3jPytwSpRklYEpBnX/PGaq62/XqE
syK5SfjYR4F1u6UeAPIDahOsmvMATQqRMPw9pAG9/nBfNO4TBpIEx2IdUg5PM2wN
+EMDCyrp+dK055RLCWQFnE6EjrXTJg8cZI27UacaHTIBupKvx21zzSEYWTegZrfY
ZEF0p6FsUfpgrBb5Zh/798YXz0FTjcaadIZ4+zZtVxlto7QOPVBpETjLhtGihJFp
k6hO2G4rj16wo69CEM3SlDh7vPA4Oz82R89pCn1jR0f3P0ch7p0Bx0ncNW6FCNMk
vrLLJbygQjyD4kBSjnmPO7tdwaVXQJRkd7CWgCKc4H0iZMilg6eDoy5x6IAauT5G
M8ydiP+LA1HX9WaPVyyy8mzWDjrALb/lm+nFYU4QApPXShH8AWyS9AH3ARBaWZFw
LKnizTynf1lbYVawa62c6eyJS8CnoS9FC0NkXMDUYWfOs+EFRUxsw1ZTTwM6MHGa
DJ1ALFT4vOtyTLqzbh+VkqUnj0KOnqDBr3grslBCu/QEtFZ2UBvvclT21ValsR8T
ta77mwtvd+tB48ECIV0msiFBTOPUXtElYje+vuo7MakaqPgTS1hmOBYmfcXIFUjY
Xu5WMPyCr1xvvZ1v7ZbAbHBO2BYQIw0WMByXVv5EuM9hW/k8axMl/dQDgoOFd2up
RhiwY2URH5iYKKSAMBypaxT1IoDFxzkFZKdcyxslhe4TmV/W9Y/rCioDr7sEy8wT
IwMqHN+6bSdjJ8auDhGjNTyowzt+v4zj73ZMdlZ4fNcVd1265xXHuHob7ngx0V4q
IKwohPgAQXjU+cTMwhGYoGBsvKF3VXL3xugJk/rQdLxU3G5xzLb44xONx9k6kfOL
9Yb3/mzpPzKMiPKWEpNg7tm1MkZMjoPwmiKNTCUpJvUxiylu353kypCEa9fyVSfJ
KdH1dRDRs7tKmxLtngdMKZt/z6SVuhn5NriFN+RnNaB0tJPNO+xnEdqK6RCTkoBj
J806vwbGHnjf0ERygcFyVkoxhYCTyrnfWBJIskDiRvcmTR4hjkH9tDG9DiYyWngb
z3R1kAbPW0mo5XRiBN2U8hIKjr+diLnRYDFWpIDGywN4zkCCnyxkxaj74JvTBo5s
bV/xUpFGwoBdRIiYH6H+YKgxEU48Wa/wPVrVQuLmERGPYXJtP93rs05fX/twVZJa
whU2MTNfi4Qt12C5mPPQkuEmjJlK9+Helr7goiESfu9/Km+C/GMrm/oZYbYhtSUW
bOCxfHR4yX50la3ugT/hRAP/hykCtyDUeIFI2sHzwss/okAbiVrADt1qOhettvyv
uyqJY50bTsq7rO5McBOGm1gAIaLPdiR8Dj1pVnQ0xewT2TMcSy7s5du87Nig7lyN
Z7mqts8snpwiLAxHpBR/O3rHxmnNp7PCsnfJuaU1FQ2xwhGIdNOoxAUho1ffs1+f
OZP7hhWFOesx6aM8WqDGL4SU8NRu2gTTl/ewVAKFTwS+uYUDDSCDuMELH+FuHzn4
tN62zrzNvZd4LEZqxZ+aJ0/HHsI6WwIc4gj26TU7Rp3+YcQQOjH6jLFCxX1Ci5zK
3W5NTnqewT+1vXO5Qnrs01AbhkltyBuua/W25+MVQqBB9UhWpPf7Z51G/t01CRYw
j3ZTs+ThfD8UdqG8ZkhpotQyNN2IAdOkLXaE5zA36m/j11DAjJghUPUYBTon20lQ
fneZB2mESDkQJQBiwi752xhr2PgJcnDE1Rx9zmPpDm8umx0oM1TqIF5GuKSIntgb
JQ/4VXzAz97lO9VPXk8Q3wsAiy0Q/36BRCQQvxSlwSCwYiWTw1zmplIXCV1KezFm
wz9K26V1m4qayxIPIVO+mVi3qQnNg4KV+sUiJJP15IkWlIVFcS0hfAkCKf50kOn/
mSmmmpEU2zzHDGAbC5CNo0Reqn6X0BB/UaGhJSvqtRc2UsscGOpJU8Gd7R1CJK+O
bVeYsWhCNxwuHmhLOB/cHKnZyJEdE1GFP35UPdDXmy25ISIf8evg2XuSCuSkj8pG
hm7Yf/0/hjNWanW56K0xQrJI/5iJCuqtcpcLRXysfxWC3YxrIm/yR5wUqCEU+iir
Nt+EIkXiIETPmRtP7JQUrYRZ/7dW3d8ELVaRnD70wShfcyHh1vc/6lGmC+vxskf7
89PxnKCQmZ9+iixieMgvZcpD2jAQ+y9mkrXp92oMom0DF/P5xh3nbwKgkS5ALtfE
dC4uTZMQV3VlQxo+H/MA4jQGt7pGKWcpHW/douME4saXmrIrm8sRUf0aXM0Ueg2I
mSQRRVpNuLSYT87qfrccGPjRcFdMirasiDogm5iPTPC2YmupMzAepkgw9NxMIuGR
4O8QpKBES29Z5xuGaqwGgc8KxhzgX5Ln5ETXf6gpFffrVes+2Qkk+8I5PAvxE/Hf
msZucJhA6qOKyOLsZvcrTQ+Hv0pFQVLSq49tuT1sfLyTHlJBpf39e2MJKBT1lSvB
qHVcaF6kdckOyjToMdM9qda1kqCBSEnJsSTiW5+pN0oR9a1iJSvFedMge95PVvna
ETfBaF4u8ANm1A7hMGymvQYKw+/YxHskXadqLALpATQxkybyWVCjKa71ZLpydWhR
CYyLxKEIzu6bn8cAgZv9i44Khz93rf0wvSIW7mTX81ufngspLkFvH1SOW9Ifgwff
EfW+mGXXeAUktOpXK8EMT2533cbluACXnmehFPEZLGEb+2ES7/MKzM3w+hBaOpr1
NBGebOwvvJQ3bkNrphr+4XFULCrM7fd6hxsXIDEJ5gmO6pBB4MbXcm32pzeBiBAE
EAHnozDGFjRWsJlQDLpDKaT0CERfEO4CgMZdirz3O0Jzb6aUuD5LyAevyybXIBXs
CtsvSH4LoVDhZ7+B8vzNx7ZsEYr/k/wdjrMA3ZOYuMKzsuXc5eyRwN/PPud7T0IJ
0tpibxn0RO8dYhj1eYhJcKMke3mBGR42Ogu3IyRe0SSvA8QmrHKixn5WG2gFMSf7
YoL90umajtSAHSR7S/trodb7iEDgWFCKI1Z42NGzLDbN6WYoE313c7Abrz6R7STB
8ZXVvrnYhreezspgcHWH6cnCeSJBYxzWcTt3MGMaTHqnkuRnPbaUwSqkN7ut2u7J
HqeYxHcV/7Hqdt81w+CCjmTUeTKfKWrlcT4/lVklZy//KO0M4uLiroS/h9s7V3zd
9gT9HfAgvyq+ZMasem3GLjTK8VBj0iO4hjaf5vS+pVuM2LXIwffRjLNjAtNMlfUN
+InJsA9sEIwaOJk896ODtXBrCZaVmWbVu8SSyLhUGBhcr3tLBbTuEFurQMTIzM4L
pVu19gdCgvNG2uuehIoy/SGIWUMCBGpAujJLS6w7MUdhsgCRnIc0zP09qEm0WhD1
deiLWlXH7zayHF475VaSxeeFSzvUS1gYuY38Ynqwu1mNH4sx+Ctxm9OD/JRBRs/U
MkUxEigUiNjWteZhpM0cUhZJxXz/ozONQ5opT/r8IRQ41gmDmZ/Pfq3Wd2xCTs6N
8nAgWk6P3kB0pdttPihK0FzugwtjgQQGQMGpqDvouLAcQtRRZIxBJBkkZwXpgVO2
HUQ19si6/lCkL6GojiAEvKQA3ppyIhznl8t9lj4uCGARvTFrrzl8qizOpJnxDKze
iN1QXiPXXZwGNEe2Fqdu1mlzYcUQo7+bkFYYixGWZDf65PJlsT/AVoZucZTwiHJA
TPmoPRMqT4EBM33zOF6qVFxxDgY/8pfg2valjJHJK38iDcLKixz7zV0y5AjveVwz
kburNbeGl+Yq5qDLuZ753dUpZzNPj/eoMKQUy0vKhZHfS6SLYDn1w3MJjZqoJqKK
o6xNZJ84REFgBu91RYm3vwHW5ClWrfrgyNK8Gl0CbTz9rmvJZPsM6HNsNaS3DXjb
I4dZFgeWbBSTuKQPEYE2E2R3F1nZIDGgQQYLmbJ0BQ4pxIQErYWRODHUD9YPpJKY
X1Nr3kvGZPGG8q9/BdEHvZeGYtylepCCGHMWVlhEE9gTqL/x0uvI7CdSpke5O4sZ
RCD671Jfdqa7/3P0gesjj45mg2boNDIPR4rhtw1MhRDjiyWp0hzbwMWAeZitblvR
FxiyxE6PArbrlgToRG69RW+3BnKd6XW4V1SqF6vwFoSBa2x5Z8ZM3mSFQYoNAQoF
eJ6MHKuuCHnlescDYfIvzq+D98DaLuHa/KRmyVaEwqwJKTAKn4xKUdciy1IJcWeE
HR8V0hOOcYV/slk6UP1gRA3bpGbZ93oWETgUO1oMbN+4PBnXGDoR0Rlan+q/RgOA
adghJz+4LOtn/cPz9/o9nYqXLU9SpaNs+AMX3geAUKjX281X+LF3gFwPQ5NZSF+x
A60pxo8kK74ZxjhwyNewRepJK/387/bORt0hNwkU0Hw3pYdZdMRvLUWSE1VlJ3Co
sb/LM++8NZkQJhiXjAq7m2ob6J8s4hNfObaAZywAwbBopx0QbohC8xbbjTzGMnpq
d4lcAugiCDhwMaSqG+hzV9E3vEOHxA34c6H9p3KiWLIDkOIKhvV84F8koPKhnFMY
xHTCvZoTE6Abp6cpEHF5iY0icjpQcFtPgnimtoU3xI6Z+CPH3x9+N+HT5jQUdGSz
ACN5sTvdYSFwCu7WrnUH5bKYQGb82NZN4fOAlLVLsPtpxUHHwvMa7QwAodV+vop3
RIugVmbZmL+71T8CshiTDO1AlQ4eDF3c3WHnPzEz3ztXlzj8tWhS362qpbe/YCTM
PSRxuawUhAWGs2OgGlFjQ5phXATbF7xgXwG+y3we4eOxo+6q/UwYlbvuE1UXX+AD
D36ifjGSs0j3Sdsl5BibvCyJbEBd49dF5cAvZLFFa3ieEvMNqdfjYxABbh92337O
wdV6//t40Z7GKhCBRsRhxgn+VvkxeYwB6lmP+5Y55B5tIBy+zqgupiG8cW4yDtuw
srfFVB9hXR7j8Q8mseSi0o+Lvc9Mm5Li5zk/tnbuS8ijQbBeJUSe9TFrhLbkS5Yp
Tzo5kNhXLK0+vGzIfYmW2aSboaERAzCadHUdZKZctXH929KDl46eCv+LnG3rShlu
I6Sxe88LwFjGsZiD4g9Bsg+TP8hd6m1j80daSplc9oO0wuETfO0/ep69prB/Oqoc
VvJbwUzQI0JC9PHLT0OHU0a93ycyqHVOWpq1ecSQrVkl4ubtZ0Kj42A3DkT+VImA
INnLM1cCkNT850UTGeIbauV+kX8c4KqRk3hPMuWtiwpb4do5Wpwx1hB2Sh4NYQ8F
bCnprDbLtyreyKBTVni0WAwtqTRWnzyzzXwXjn+HRXl17Fxu3Xj5i/SzR84nuThn
he3AhAQeOXnALYeC1cq0kc7YP6yTt2PtvrAN/8w6y5slv163pOI8D6UTOf5SYUMD
Y/WiCeW4JzGWQ4Au9XqX5vw5/0th4m4AmFQ86KbRXSiRnMS0n55XsKSFIxqXZTHa
JJknUYGEAfLH0MuNNEkzwteMiNXJaPmTrEZPgL5h9G42sF/LwdUgkcLrNCqDtD8h
ffMLLUzdMJ94WYoxW94kg+AgohzHyvAckZCEu3EU2Ei1ds78CQF8Aq3ICQF1eM0i
BIBH6ZkuLeQrXitTEwj+hyUKoaDPCszEmIPFfispSmEMhI317MeNJ4Ei1jAeyv82
R3+vfdY75gl/Mf/I6Cj6Wc3Cj+S0UNr6aA3uxE1hd+5TBujNEtwqZDlr92edbStc
Ju841SBljx2ZZF/MKx36fMWSa6Gyo7AOg2++EufhSzr+oiSjAVwcieCwms3qky8A
T5jbV5EF5jR4MSJv3l0lFH2iK6jlxCjjsPBM2qBXfSEPURK4mxKrFfZ8yHoGRKsg
ZvYIx+X64PiHrKBK2p/Yfw0IQ1wmB+nHpJjrP/880/qeSbgvbEOdrOFbQtmmxhEp
+vvmNz8LwfNHXMsqHBbol0bvCCWBSQdvP6BXrMnAlb8jg/18jP0aMXiOBiXmxNZa
wjiT70HitLJLvplLWFa4dGnEIqGOxSfk5JE8agO7PSGkDpaq71CvLiDzMuMHLMo4
2L8KnXw4xKql7HMzfZ8PdbkWAuQ3RhTJsz+xIl6eW7f16U17/xxtB4QEMBgFBnvJ
26XX4pSD0h8Q1TrOty5K/CptDVT6Z44UsQbMMU6+RSMRf3+93QMFajkAZxrYlddz
EB22/y1utvYJGiMLqjl+pNHq0szDfHSPISu8XkjSC8Bo74EX6Zovk7Jn4PIYOAOS
lZTcWgOboSH3PF6NLC79RFOSdHSubRUrB1/kdPnFO3jnw3b2ER1MX8RL1Utt2cT+
LgCQkiYbolm3aI1TRRWkXBpp6Rwk6OlzhoOgFlQsktHNIfBiXyCgonABK5B2VQyb
2B4twst56yQQCP7t/aU9EasG3GHdWYyQPDkG4yX4uvyZ+4xl3ZXA2F/nNV8Ntz8P
ldqYtN4qQIfECkLcJhAkA0CRLcmsjou4ZAUUylBhrvbPWO4aTou4+SKGBvPzP3Qh
bKuzMYGx1Vo/DQTe+PWznzLDpQj84ZWpvVz7VtcL9gl8AJ4icgp7LiwCoNhtl/VL
GVJDAlW1CjHlONaj0W5qfcwu+mey8+5gzaBBGEnGTc4/qegH0L1sFHDhFPG9MI6V
wxv4KMv1jLnhST52UWmme4UYZPfvuJigI4d8SWJXHWUoRboKmF76P7IKEaIWcBbn
H2IPqRk5wklO7lmtNWVraZfkl0x5XLJhbm1a8tKWBeGToeLkFVq11FFLOArjkCSU
RgTJr5dCVTHlE5sJAcF2GaOit9AYsbeDS4VvXf6lUnRVPSByyxRfC3rP9+VsLNvH
JZvCvYrt5vgH++a8ji+4YhsoGX0fGJDsBqeoGwN0fheY7ZL8uZyGyjQNx8FO/kis
hPN1+x7RLsooA3i0VaRMjAePrg01INyW66gg5d8ydSQavxShwNnmWijEQxDsq5iG
QeF1D7UHAE3VFxYuFWr+rQ==
`pragma protect end_protected
