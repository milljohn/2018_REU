// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
X5hU3u95tW25w/NvvLWKGc1DJ/jwA/7MoEPygFw5efXFXjtQ1GRkCwrMxm98fd5Bt4DXQtXO3Tju
ec6X2AzFpVLyIFdYcelXaqM7CJz5Z472RtqN1UXMEwtsrDilb2Cjms3aqbW5azB6ZWjqC9eERhfk
1Gtb1afLF6/XcJqiqzd1y1NGaASKV4kxgRJrIMFGochGmmrAZPNBaSKZ3g2hsX92aMmzK0IujdcM
d0csABNxCVdm9NTo0g0MO39wr4JOyEQyeVyIukZYMNoG3iWU4uC8OD4jb58LWnwPRIPE+xsI6yYi
AmUuyDcvbnavmO2No/yKYqnWNsO+6cMnh+Qxuw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
T9np9P708Ee+yibQS6oVq3OdY6yA8X65lKt4LxrxFBkDtRJYdu3R2wqquyjshOw/pM6Oyte8oZIk
5/5hT2AcFs0GOr9DfLIeLDEwldiu/2mNLiJXAItg488GC09CjvmDBD1jUQpRYYkzmL8O5yZorjEq
QOSf7VZ3hshilvpWcoWYFSuM7Et+Bwu3k+KdcHqI/ylNl2MUm9dDFvkT3/T5BC915uKcnh8wOAfM
momA7BGr2jss2FarW5Fv9ZdigxxagA+Rz9B9H8d7dNyLV/350DVAqayEXoHq7N5L4AbnM8donTLc
B4HtomNuLFQxwGuoRD8TCGsL/NI+Ddl7QdCxwEjmW/Ylg+It+qIGnGeONJvlFt9FQ4PUAbxZo1Ca
wmnBbU9Tn1x5oYB06d4dIrIbzmC/yo01CbO9olKqAYbqeGUsM4oqNs/AVRXCaE47muWlj03AF24Z
SYhrD1kDBkrhwk6KTIt7OZgZRr3JjTzYxqlZrOlo8wxrq70+1qlteyuAM6WCaKJAWXKQ3IxFJhZp
sPiZ99oMeVUThPE8oWeHoaUqD2urOfGqVJg85IEDLRvf94eRJjYJcO1D5b8s0YMkgUKx5MdgjJw+
AfNVvz/++MApXmQzHiJJSICBxrzLEfyw02UpLu9d0WUYRje++JSP3bQWhMqJUTfd6HugTnEJI2vv
dFx0P0JzrRhp0AjwGRvUzMtko+LugwfW1tDqSvx2Mr4PgdYHpcGer+OjpPTPjbmzlGKx9SxR20S2
KYjYh7bwA8yRqAIajOvNgLBJy4xaoGIzWMJ9SqzD03xXWlQkswTFDU5iJJjd7jtd1UzZfm0O9m2p
ehlLiUovPyyYKR7LUDjtfNKaq72r4TQ9gNfv7wJ+upzsccjUZi3gfbhhNu3C2TG1UMThmk2Ab1Kf
Ugf8+tMtA8dZWC52OkWD0+9nrkAuXpCxgY1PODkDRnOKIwSea/mUk4Ci9fzgzSSWpzhfU9EilmNK
jCIdibI+fpK8nKafyd7PwJU0wGp41K1TIitJ2WiaRWIQD91XH6wqLgJciLb+mp/h01nWIDrRMbcJ
AR/7aUzVDXYsP2Tu9wY9oKGhxrMrqUMtuspPNmkmKwMpqF0tj/A+ard53uh4Jgda5CKgUW7wA8hB
O7TFIXxwfaY8QoGN1V3F2j8/dRWFQ3jgM07EbLja9t/GshRE+YserZqIMjY2wCWjVb+U5t7NEi/K
YJ6LcEYJD2ETbJeb2noiLk5ugvbR8ZgJsIxJvJhnOG0zyrkFg1zoPFLpTeX289c+zXcwoS/lzg2I
fePyjEi6rJaScCU2+tyBIM2ZabPTRBO/gTQtsoxtxQZ5oXEbTPaCAuVbn2YX8legv/125gcjaM18
USGtsOaZCpDwrPL9rbjD+Jmq8u+B80i4+C8dz946O7iLLFcektT2Igh5b4/5tDsGqOATqgm0yeTt
lpT2ROsbwoP/8oP1E4tSAJh5j8KfjOxvaSrm5g3b16jA0JfWrqihyw+9iRnPHnhft1/+y5z5onTQ
1RZOaEJ/1kwYz7Q5+ulQHWKe6KeQScURIGLjzZQ6LhkaD2dXEe8SFoFoz56c+WEQ8JrPB9Ls23Us
dir7uuVJYckJtnKI5JesO5FApQL4X7jkvj9IcEUk+r3I4hRHNcT+BqeN6lcKMhBwoO0RiBA5/VxW
kW412MimQM0oiHidqw5mr4QSPE8QghYwBS+GuBDhIKs0cG7vznfsXlVZ4rU8K3CDQspVcQ7Sv+Sa
kPNhpDg0v5oF5+Q/+XLrpUaKR2xUhLZigEpb21/Mxb54GwTqZmVZViz312bR2tvrOmerTA8LGoUo
MkLWvUXgw06Id6soR76In6N6Dn8AXw9yDHvGiKRf6PIFE1hNLvOCX5ddp8p82EQiNjqMR75Qx5m/
1B5vQmjtPHZPVCXxvJcU7DExxNJ+kQ9+zzNxmPK/tLe2Iv4p/oSKYd2irjUOIqlJ7Vj9bBvJjmDZ
rd0z5nRWqc4b+9MvPMDxXbgMEcQw+hpj6mTLfVcCzXg5oiO/CPAJ94oXc3Oto/UxWExwvfTPvLIf
TdhkpJO9vEUz+OvMhShqpA3M1PogN7G3aYn4hmgQQv+zbeDFmuVL/O+rZBS8qKmpJN0k14kYtTYw
ZioooFZbZ2h8o40p6RDlPdWD6kONYQRoTlcaZ2woijxQ6LYloaMXygLZLvbvqO3kdy3sWIsfKAc8
Tf4J+1EM+0S8CRF/tn8EMhczeRDjRIjakwr/ZrbnL1dbc8hhhqTMd2UoIXZBNpEQdSwy6tc9GU/D
rCtknUT52fpCUEOxlctL4UyTykfQ6QhBoP0WdJq53g4kjhSxzuthA/LZp7BkFtte9nPUvtO5cMV5
fK9dDJGvb1gN4esq9TBE0OrlmO/HaA0cnx0jSItOksx9FGk1Y+ccvB7c+0Gp3hwD46zhT8YQGq3b
cNIOFqP244L7VaZkY/txdp6vFSNz95/jFPcDLtQZ9cpFZtDbyLvG6ZQvqAnqTL1fZx7LSwFJbZ37
N/Ej0p8if7DnbdM5LonTQpzqXYd2ApuaDwh4DiQbEHMmEoR/1Dnnhc5dgjDjw8H9VdkXRqMA181a
T8BtW8QZdr0DpsbPsMooMS8rC3fzH9oNvrSIIPavzKu2bNJK9qCxw8hVkugWgmci5TKDUBfygRAf
x1I+qXst21YlcSbyRHkxJ6Nwdq4vm/x2UAcQEVvJKG//61TUtLC4lT9lM48YvI1lRv1LyWd9mrTp
zkWNNffQzlTSjUtsshtRSFnCmF2UF3oUKZsYOU5/SqZv7Kc6yBZ/IbCqqpg8A5ImIDSxWyizYsG9
U4Msed1veYYQnwBRiHCN7NnJ4W/Ku7uQD7PsoKxMTjiOEGj1bdRIA+Tdd2fxon3WHVyZdhusrdD9
LtvTbOy8qRyM7wa7lN/JFRKEZ0UzB4XT7gEp+rKHwI0mUj+CljilxGgU0WVqblgcO5iuMOpH5T8X
ttK99mfSnsImYYGK4IbFu2DGT6qhBMwSbpsd61dQBarHbGyFTlxkAahO9PVEimbO/HbzoZ8CPM+W
UmGn290ZBeaYUxseZFKkD0eUvKV0148c260581KvgIda4sOU8m/DYCj3GVsotw1eY9Gp1sNNoX/R
prUECYpMEZ7m+ja8HVPLSyJG4DT0TP3iauEDubvpVxldR2QVs+WF+5qN6Pf4RuYB60eFOeaXAfyN
fW8jbNn+fMJ17oJIvSHd5WNEuUV9geqIOhuZ417YWTk6Ff8ZDv96o6rV/nmE5BFkKAFA4ermh51A
9ddWCzW9wgoWC+mxJ4LK07kV+mQZ797dVVZbFpm1c+Hg8FzUewp7YHUkMvg9T3R/63McqAwhzJW+
H5C/+NyjkiCoUUeCIzMv3wbl+i9S+Ug8DLRdTtmU1MITUJOl7gU5QueWHKVuMgQepNLbo6zdMgw+
s84Gu24sJFcvZqX/8exoqGMLvMQep7a2WAJc57ulgb4z18zC1VT+e4Xe41euFAK2xH2j8lRAod9R
Vw4qWWSDJE5GGV37n5lAj61PDrcyQEIiZUD5T7pZMJXjD/buAcvresFcYNAiBkj57xEemidBdmy2
WdYHE6fHQ4Z8jjWhYAvqrQeQIHBuy41tnH8XRVFTGw/SEQIhsHMfKzDe0bz8sWo+uM5lVZT73Jym
ZZSfBlEZ7+W67/wutIzNyOtg3/cAoKR3ihPtmbDEn/E4T4fO2mvg9rpgT7FVPaFEC4ANt1lgZz7q
R22Pxoa5JzEfwAN/NltsljER48nZlZ2FUbv22a4O9leVeZgSb/hl++JQt/Qwd964ScltyKN8y83w
pV/62E4G02626YIjex29VlaP9QuEfVbxcPwv/7uWK4Bc+rAECKuThuu+KUAqi5/AaiFfrUaBct/L
yVt9DmBY338heaOUBs90t16PPt2NustCf7eLCsEJQjY/ntJ/BaN+IbbeI/sR9SaRteiiIkfgbbW0
Mh1p5c/h4sbJEB7d49MQC7xxrKWzVTJp5w3l7w6YTnI38Glhf4fT4/cmNejjgvfxfFdeu+r+3lRh
HkuvqS0jkARFkZ0Cserq8hTBI7LaWuMBsgT9QOFmGSoQ9B0Ad4HCDuSi2kY0dikjp8c6B60B3378
TIN2qUsx4CzLSJUfBph4rJc2YBDSOADUhRmTVtahx6ydXRPFfZW6GxtPxXt+qveaHo+VSAbMHCCw
MLGh4dW9Y1WD6mlMh52Y7toUpHxcaqi/0FXKDCeT72r9Mfp8EoWkF1HVz9xeWfD8s4eNUJTcf1ex
trSFlyaO/N/sSrYelMf9B0F3zTFXXMSYugmGmv+dD18VHTybrG69kJiurhZ3nydDRbzSaoj+Utcr
78MufaOnSSkm8PYPMh2EnI3M9/JwSZzxKXvHAly/SoI1ZuCRHFz8ROu04gYCkxbMA1eaoqpGv07/
b1eal8IhqcPWuIOdEoTP/YFSPSuhMsUITIvN9u09FYRnE3QMsSIKv1MrrZJLum/BKjkTVHmtNaQC
6NU5AQc1px9Ua660efOL7x1YLJenkFk8g1ogcbeKUI03yOM7r0e/kikkdGeEo75zETc7tU8azXiI
/DmZlZA20F1WaksCMx7tIcnzuUKIgC74lVEHk+2XPR1jP40MONQLxl+Mp3CdKfSnN8n+inkOaPiP
V7Crr6u3pRqAjedPuJpbgzstHzClvwS3/SlDARKYCn7eygzhw5Yh67LWTeA3CyjptEEpr+tKvBYU
EmjzS8ZY4b7BYkL/F3n0OD/HfieD8VMkdh9hV4oQ3Gz9P8W+6cUK43OiZ6p3/IsbT0uKoE3oxxSp
jUnn/8V2+yP5tMDFIWCI6+llWXKreQ56y2fwrZZWFzlWzB10QDAiOkt/aQdl6lsYwWYl5aYnvUlX
EmO+9V5IoLZEli82JUUsW7DzjjE6IqtE020g0luUw1vC8yzBpOrhExsUgHpI+saX+2on0pGbICHC
lstUg0NKAV17ghwpkw9iZnBbnT+cPym0j6tEYzCe0gnWLWjmEh1G0sQm9qnJbwVMiM9bZ2gpXTrF
iUl6675O8amjmMvZrtNZWer1VnvPUBOP50yPNR3HQuoPlzbSvHV/b4QNwaGY4p8bTG+T0NIkyrN+
aLbHPh3AgMph5pTea/NCXtVxLDkkcqvPBwupkBvaAz8rw/no+GPd7t6+UH4vL8YvWedm0LUQbm8Z
UrgEwsXoEufTQYq2ebBhhwfdyL0fmsNHoPo/Rd7EfOeW5R5+PJnBZ7PJSx4azUDiS56Rzdw/HViX
+QQX84yjexNKbTooHXb0oa1rJGuvdj79Nn7FkDJqod7RIPuqWR5uFn1xxY1EwgR5u0g4JjZc75R+
u6QFKG3T+ILNX+Ff3Aylpg74lXyf1LzmrfCI8GDC1LaVRNx/+IoAliLkPS55r+PygeIqe0PeqMsN
n4KGRS31FmZ22H4aw3n2wDc7KfZhTq1l7CMxujUJEJEt6ZDcSDOiEqbNVv0aCEhC7TIfYCevJQtO
RgThhWFnW2srzu2I5kXVGL4hCLCXuMG2YuUIgm5XyUTZfYZTL4Z2nTgwqf99A7peT160yWCeuBMa
bWk85/p0mcUDumDcktn/ycYmJnO1T5jci7EGClgFfBX+E153529ZgVseOE1n3zEXtb+v92UjN8kM
fktuqQCLcF5L/iFxuMBQa/xSwfoRSb52dp2Yel2DQKYFTkGVpJ4G8RH0hlPz/8DxvdClmcA0TVOD
IR8rBF/V2zLso14lSzK+hq+3+JDAGx1J/xBiJp5ebFVRB6QK66S/y8PfRYIotG8o+GDCKwe2rUvv
abISj/q3ts74O5TJ2MkdLh/iNXhCx7nnI7DZO4EBD4/BEIgU3m7nuImpLQBqKWxoIDZzed9ZGllX
YrMWmAfTZy3RoKr1SQ+8o8tfJKjLssstiO5FJoxs+l5zovYktLnbTlKJ9XGUgRXJ4bq3Mj8T4J/T
M6WpCwmFZq0fRute6aF/WVIoE+upfTc9YxpfotYGG7XobmVV3zYmPocRsE9BrTQN/IlgfZzmZCQy
n4m16p2Yt44WhPJeHfcHb7XS2U/ogF29tHfjh/kVjBT2RQvq2Jf3H86l6Vw7+OOvt/XVZi0wg2jz
WOGsuY+0E6/95nYUAi1Y6Mi13cVJuGIoB40O2kXO1ClazRo6iGi/19lH9dMN+/75ixiuI44iyf20
aykeiv9CQMFRCx4EGSvDMeC9pq8dQvfBsRnPwsFpJYSUx0VgaVwS/BUDB22taRUOFmEbcgcJPeiw
2FL875HVB4XLydfEgp/pdi4yteng9Gy6XGKoJh8Envt9x5sQWUJ4qLPhLGH24RMasfLvq7/YsKPm
9VnJrJX/AlwHescHjBVjZlOvSjs+YYal7v436r+XHQeFEMlr2LTNjBCHhYQJRYSihzPcHZDA4SV6
7oKdV51EbPrFUUJ2eDq74Fl/DPiiIhsUvupjYaddOuL6gwZ5fTC7gmkfVfTG5c2HisAY3h2gKezZ
dqHkpM/IES9S5m+fw46lfFWOdkqPEC77JQ5AmpNgEqiVHMBH0T/48QfQ16ua/j/uRi6NT7XNgx9y
UZAdaedlXD/wuH/oibyzj5sX9MUyWP/kFQPYhMIRTxK7M3gJjEg6NyXbkDXP2+iGW78Br7flThad
dNXUmqkXuSBiDvL6g1rY5Eeyx/9zujdpqXfne4Gue5QAmJnSONMUgtrcd09Ag3pw7MuoQEoSTG/P
sqdv7SvgJfhmZkCkit4OxDL6zWrJN7Gn3ahECISTFC5VLlsOEuhDrM0U0vS/HGkaOKX2ejIB9VNH
7SBzL0q0TaBh1wwtpV2X1R9ahqXSH00w4ZSEnANS1JvgyM/odeglTHE+eKu4jn5b04lv/wlj9R/h
AULd4hw8kMLiQwFzx0Ldu+6aaVmk+I3GpYLMo60D0BTuhHsdMUTF7wN8uxJA1QxV2Yr6zP84E5OJ
kUESldB7Wmy4BJQvXVjOyWCffoqBVJlN/gZzjCN67Y+xPXvtIXhb8REZID9JtYszg4LddCaNcCwD
DzIzHmhfTSJ5aC3okWGHwhfhjlkcem01wkwHRxh/YWNRz0wkjqVT8hKKK23uWDHbPke7yqxw0mfV
nw+wMF8bEaPMFg/pk7v1oI3ALZBJn+74BLzcyQRW58nrkl3wOloUyivFL62ssTTehQEObsTuoLiZ
zmbyfwmUmWNYck9lGLW0OrEfMzHo/92rl7+PBHoO8Zvbj6y94sN2/e6OwpQnjbbmolF4NzT+/PcM
yo76pgqhdtZDg+nso08Ms2LUB3tzioRAzJrFb1ZnHiuxse7UiC6u6C7zVqhDS+hZg22STtdZp9DD
0ShlxoQ0DnHRLD2dFmTLPoOAWwSq0KJn6+t++klQLxx1XAe3Fsl3SnYrC1eZG1PrUKN4l4gW5+TN
Ry18vQaCvBcjyl5fTFEmrga9noPfkpKFLqId0oreHLWYIC6sWWEbqLUIKlsyyvOXBRo5pSAu2g45
qdE+1L06aL/WU88eL450xDlIsurqlPEloWo9Vi5SoDJnyUMKEhwGWaGQebz9ewOk9vvOZtK7kPSv
Gt+7CuBshY+m0vMISlezL75wESTnmQdHRinG5KGZ6z+ZhJ59AJORcEm6fKzdqrlKCt7vAT8WNY79
rknxwzalTEmf5xd8Fe4khXr3R/HTLhQ0U8jUC5ROGKfDACO0vElUkk2ES1egTMx62H/oY5h4f3Rk
28oXNfHDHlSuLmd9KuobWmhz/eWZajpEH8l/Yv2ZAyKQFLFpHJgtDP0KBdqhYiddFAKo3bd6kewy
t2vMlJK3IMSRrs/JcXF5+pphac5I6XqdIJWl8mPh2GHQTLYdLfAHwKNffdjiR8t9wp+LvsqACJ3P
VvY4It2VJVqGoWljagckpaFG9auSLJNg1G+7pXmxQ2R/kOVSSlXHUlYutb97Xp8pfYmZzs+/2PYM
54HUzU5k87nXqsFtsgI1vgfY9tc1qAjehoFKh7YMyyvxOnLzuQ0eHLoaCIg+9JQxlVThfkKTShsh
Io+8O9f3Tlrvp0n15A+LZaI3uxJfpawmUBaco3xE2oQOeJhLNpE33MGviIgBVAuGEPeSxE6o1TVg
cf1+wAsyuRyWz03m+khsFdpWZaMz6vzeE4sRyPem0LoqSR7urVDm78QgWYV0hBe71RhTplsJUJsv
qt2G17C2oD6uuIVaTu6Wv92syqzw3L031fR+gXMV5b4beIRwjTq1j36eMCJrT5jXCMYWhU1cjiLb
oO6E3e3iFGZxkhSqn0AH+n6O9CmViuMrSRlWv41hGJzJACKNQ7sx4nTMMWyYIZd5Iy1tMo9uVuPD
mEd6mqAmaPZuFy4qntD3Rmj7333GrxVp5UrKUPwhsNi7nOboeqbdoSsck6QrpNDQXdBd+eYrDTht
nnDHQdtclD8Q26PemoCtEeFBUICIRIREVmD3g07FRwuUTUOPJQmpmlRSq9lLkHNsEABDCYMzbPgV
rQ5jH8M0JGMtbb4MS5Sv/rIlpMc4bvgc64btEivo4xdRLtTOCSOL3dA2mLK5yky0l4KTNmd8y6C1
ne6P+PQ8uxB4eEFFcSFqDNG5spKSNfXgOKwCn/jcPEFX7HvFOd5EO5AdrJcUjGLHOGK4k6yXGdCm
CEayLmHbxcc04rAjL2Y08HcxtMom/CqO+SCKi4wlzA0+5fMYn4YphF8/7bR0D/KYCcOUdMHrTeWM
TI2Os6ovqxt/NN0c4GuKL/W3bmOkLiDWyxA8VdgivX0cjFwiQNx5AEDkheo2rpPjcqEXqbk564t8
a8Ubumhr06mhkphUamTvCcTfVPYt5q0rFhAYTO8T1vDULNTdk4L1sBGZ7vWQA7kbEOgWgEVuXHKQ
ESEkoON67MAllLOAVMNzC6+O8DY5lzPz+tStv4fD7WfNp02FDV2loqjvuyL1ghMYZUNGWTi1QTOL
ZVaPl78xJlkElc1STW5aMRmtBlz89REeVAEXuRJ89xOOjlZazlWdxKKswxUnjdLeE9rc8d9CIkgX
MpMDtNR3LsEpY+5mwUe/T8mbIGWlFmVjvy7hmcqMCiBNT0MuoX9XUcm9OJFXuBr9AX6X5W8swxax
BzbPcsUyWDci+uCgcvQGFrfAo9MZBIlAIjVlhzBJUKB7zg7H1bnqr9Xc+sSPeja+lnS0LxfFWnNW
N3ku8zLthb92hXDnX4gCGVR9Shnqm+dZ3HpGm48TZ/VM09AYET812JGlohfVwu3EvRjRjCuNr4aw
b0kGp9iIo8UVj0s2d1rpJrI/a5ks1AMNaGoflIvKL51jbZ1k9xzjM2o36ayNsYgCHvAQnGIcTayO
7XbvNFtTFE3jEpKr/7kYOr68wvW8j1etEbuxzcTZVyXQRpHWTqHU5uiWx5z7qqPiibS7pujdHKqV
mbGCzthqyLR/+orxLRJ3OT4iwgY0GJouigo0M0w1IZtYz5+6UbZWg137QGe5OrzgHy5JD6gEWJ4M
U/2zmuVa4ZVDoxQF9KYZl+3poLFfE54jFgwRicm0yfwHW8KFYD0AGJfB10H6z2GbA8nOQn9Vw6UR
nVdQnM5XpYn1mxuuJuppCiBtmi7cDjgneDyMVxjeihY3HpJXrUTEKrfCgogYt8ItRpCRqkKqzunq
t9+89QdIjC5ADsstla8ITsiVr9mxdGvNDyRxvTwlsDc+ALZPXnWz9XyOdcUw+VwcRJ6lDy3Hh9cQ
XGcI6Xux0t9jBXBsXKvPFlczeR3GPrsWn6ODb7KG+mI323/u6VjhU1vbPc0iUFifTZMNZ0QQHHbt
r1PZC9B6wa+714m7zne33ZB7qJbynF7K4lRrt4N6G8hlUyKUId96j7Lh8q9AQG1XinR43yXToF/E
asE4B2kSRLh9qKln3pzmBWcly8/qoiJQB0m59YDJ2hf5In0wIk0D/yiDiF1jpS7ltJ3n646Q2NoA
iWucZ7+4UDIh/fX43+UwtaAPJokC12BWiwhf3OvkF7APKDzcbL+Mrxg4SjZQ3eEpWonbAiI0CkoG
4xrulSVhebK7Q2dSVbp+nZfsaWhjcHUaqCK+hu3HGVQihOGmlywvHPnyM1ijSyuZbAx0IVe/GMQr
Hqg80VL9FAvc05GVKFFY2ABQUxKNvSIaao/21WrPM5LvwlMXz4hRjU5eYWkHxxevjbXWeoMNmjQl
MaPMFyNoS6vuyQsxfeqqckoUg+tlQ1Kx8BB4F8C3fmXAMkT4r2YaFbulsbGL/vGzdYHb0A4qbP+8
2nNZiJvuSUSoTJztke7OJVjvawRuyZ25lKBs39TAMf2Zo38p59YRpIb9wzu0V9xlb11WduHbEbpk
tkL3m4pYZrKUIvwSdZ+cs4HiOA+clE+HnxvkWQLT4ziJEu70L6DighWeHIoYxmlCRtlC916gyDWi
NC0tD4i72ThXfrtVoGRdEk6aeUYvWHQf0D9zDBKItjIi4iBGpdUK14DymJk0REQ7uZHPqIW16wpp
iX5tD14nHwsJxanBKC8w0jkm4cbybgmGX9e10BU/owRNW0tmui9B86XsBGB7rB4kn7KJrRYNWA94
D8D4gjA41MPYl0/669Z7PiI9k4H+fpzfGZGc9NKKZxBRiNvpgCN6K4X8JEEm7P9I2NjjrAvKxj7y
Usq22fioHCGRbBcc221Ik1uIKU5Viu9jZ7poOvgap4XNxjYhFsWq5rvuPN0gwkQ5mYATzbOxjvce
SYuUGdJ6ds3FLzU/ULYB4vSc1GvEK72apDN5VdL8IDr2hsfRG4PixzbmSBVFp6VacQKYN+K0o7Do
/6K9BVPuvMFZbbjkHFBu8IKKiQhAQYc7BSBZ1VZQHQF2y7WqU3W1A0FKZ/rGFHtnl7L92dzVQtLp
JUCRwiu3F3ZtBhCQqqjQUIpYPYEVTArK6dLJ2YoSx700BHuE0Ub5okuCIZ23cdbDRd/DpEC34bUT
FQP5KrVyj3nA8s+Uj6d/mIck/2mDqiyh3hC/tprjzgAMokKvWcIo2DtmMNdzWDPyWuUIUTazghhu
KeibtIsAz8Kb6HSx3idFWpRDoobkxMbb48JTeAMrirBR5Dr6nHezcr588k5OO80X138/pbquNKJ1
KNm89R7NBgV0SzFypJLmP8TsnRdzkTvo/I5/IDs6s5qHWjLf3QwxWhTx2kUT5j6QAaCpO385ZKaR
s/txNRsoKL5g3qhEldL9JnNVpuSataLLosHz8aU22RS+BmFh0EhB166UZzijXk/+pj2Qc1zcDFgt
p176rHOgmlv4yuJKiMyUsGkBXMjranVjQ5sB3djn0vsw6iPdo+R8dBvdyD2FSTZhEwcuBZJYWPJV
kE6UbTn8LPVJ8Nwi1BaGV2yk/O+MrL6t9NgRZtOCXQeTpKuKBdyaovdcHJ/Y6TJdRPQ2NNAQGrdl
TpDhb7mUYHJfsqDd+Is85FyLGnNdKW8QCIkpEw+JUYuLF8vsl2HVJxSD9jEfHMOp7Ui3Nch9Vyyc
NdI/niqJvARJp4Jof2BHQkoQuAiUUPVJ+kN7Nwp40khfFoUSwa9X+v+Cu5pUhRmhQbOPO63yVWQu
DNpjI+EBNZDwJ8I7l93UvnxFldjrcgokUuOB9hUsARjejYJNSG7adIb0DvVPAP3JrkoW47lLpm02
xjUhf93I8FqVGo/VswUU1yqleE04MDR02ISh598nM7tRWOWeGdvhn2huwa16dAXOMOn4BD7mlUPt
YRXxOFv9Le3xs/MlczL2OkUYkq4WEdI1L9B2aUbB50sfpB9wYWAyOEHmBzNdey8KcqVT/TjoTuer
86EE1J8b5/uyfY7YbTq5ZTga35C/T3GpncMsrbTT0CCOLjhWu86J10bvqnqMbAAPoIPa46A1+RRO
2Z5Whrm995BQdAB3JG5042cPvjJUeh+bZKcd99pgJm5DsQrnKvBs183gTlO4PApHmrOU18wvcHJM
wQx98lzA8hidW5+toegwzO+AZRLtZEnavKCW6BAMhtPN7Cp7AFCTds5IbRixevmHkhF89BMRzlU0
fBZrolclxVLj/8us8CNwnYHQmJEBcbw4t6EJTdpjw8/4PcyVcvaWTxY6Z7EtcMrYKFv8yVedUjb3
+Y5N81x13rXgE9zWQsj59dWFUw3XMjx5fhsIaZlaLpozz7k4sDz4A2Fxz8IlMnnrZZQnA6bz0bzl
oS5uV8ffnKPcZfiKBNolo8rkc4p4feY37WY2BWpzWz528eugCJfW7Px7twLBm9uWCZY0PhA/ZUwJ
b//c921MvoyS+6l48hSAf7aoVrE0liKMjq3VmTVbNzfpnUaNr9payJElDNrmy4WeiPmvtCLzV2Ez
TyjxY9K/0/+V4NOk/MfzMyhkcOlDzAx/3YNxuU2QDHrtp2gNNt9mpQWedIuNJYvAajAPodQkLaJT
Zbf7IpiJNlAXgXqWHCBxXagdQVdcqSIb1CkImnvKqQmmKda0DfMd2PIJd5QzTRwtXdYc471Wx0ID
7X1AyR0AgbmwFIaZ2xM7OCGx/EVu62UWWq6FyI9wMhjeNKeJmOBdo2PY7khlQZv/NvDzppmuV4wd
zVIYAfoJKc6LzPtGKyxMf1AgGhhHxzAVn8cT3t2JoDu4khGMJ0/nGdGTNTbSIt2XoKO/5BRmtcEX
/G/vUi7JNRZmlo99TYVvmsAVlSA9bD+vbCCaD8I0ZhLnOAWdeMBcr6eZ+VOZwv5QN1TvFcxHA90S
hAtNSetbckHZ5oBO/mnMrGJKQnrHwJGCDoZEPzxiJ88UjxpOAdBumILaETjyh6BcdLX6nEKXlaQb
JxY/p1Jr/4RShT/dVTLXO9Da/b62HUhGRI4H3kvzezJ+XCbKKmBm+tj3wf0MvMDJRX21yh/2yya0
XdD7EIh+F14h1brYbH5XZO8oTXTkWWjWBWIVAfnyghS2vv0CIPFySkEuPYA4RkQcLsrxO+FKG/fA
BB38TNOU9WTziPcar1NyfTJDNemAv//9nELDm/oOvMnNjbmiyRPsK5bvOxS6PjUnALXW7SrluIcS
bz5vK7PnQdXxfu19cyvucI1zmzv4QHl9fMU/HvN7kT50E2sMfyr1ppm/edwDc5JQ2ewWnqaQwdD/
04TJBI6HMnd764B89dTslFjyzqG7SN233jpvM90yhB454HRv89i2kLbK3zxM5Y9WPMqfyIN99tBw
7fvHuUKu1tnhP3hNnJicKQ5P/pWar3M4U7HNUxrXEOokguuY2me7r2XfYZBeJuKkQ1ZhlvegJy4h
m2NTxLCPpnb+uE/dvNXk6zY52NFrXrOYIgqFVM2uBgBiZd+JnCnSZa7vfqPWexUVQ/Q4NIF6aPFm
xC3IgQ35Yh+u52PEOqNwT18cROut5pXxXcgBtVjgyrrkTgVaOOILI3QrefiZubCEIaoDwEoq1dyg
SDkRW97ITJ6co8EA3+Jo88YcGUpS0DwWksqJcrdMxBOIdkW74YVFoFyTEddhf/vRTvHDtyaB8uin
VV1rUAiKX/2i/7iF/Y2iJi34NZ+vuxKxndK+yhaediqobFAdNuMyOaMGTi9bL8y3hPqT0KjSi1hf
KwTOnZJuCMZM6DHlNWZMqPVoeQtu9YPj9nALp/eE1bvv9zYqUsTFw8aZTvwvfPXFQC14FPkePemK
zsGLjs9i4xGGHSu8dhxbSmhZb9l7+HWEgXOcomCsx4LUxAiqlp0Wk+jdePXpnWygct3ItsRIutqs
mgRvU+ZAcY5jh3OXEoiAAwp6SRRPO+XM//qlQLGmTLdl1GtmU1ufDXydoWl3dbulcPd8DIIp0AJ2
BnYOoZJQJjgZ4Z/IoAFssEO4aSvpAKpI48SuP5mfk8WNSSqgW1KkO8IAmd1oOiCV0jsJDGBJP0cU
WxT6LYOKyJhcvogP4uXDizvpwoT3xdah//1RcPVzCXc09DTWsk8m6geONrMt8q6+IFqkbmgXGerH
1vyhZVBr5nOZZqcek1um8kvuSsKtda349SgFhGQXmIrtlgoCN4p+R5PJH2F3PkenpY7orUOpkMxS
Nij5pjx73r7NqBPQWmmILOxANvlYQShJXuIXu5sFT7dRfCoxnx4NhCDOyH0vKKpnFk0lWTemIBgt
eETUQTMi/G2DI8VNFcEp8oY8ZM4v29bO40K4G/EzUrCEvK29JnZT78GIRIGgOAeAq5YPwKsDUnQb
Vx9UGU5TD6WjpcOEtxpj6HAYy43lNHYwKzn+ZmHYiVAwr34Rr5E28DovdAKGnVKy97XoA+EaY6bt
xkhKrr0vqb+yix+6KKftjqC2zTXrvNaoRkscnpl4gle/aK8lUHQhjf561GXHxC3Hd9HOkC1RlLSq
6x+lfLEPxYhFsT7toAn/kANz4fhGKB+9HgFThWOj1CveMASnmGO4JeDpXRHHj07DEtFbp7C7EdDZ
JVC6f1i5+9S/BdfgCpIY+2YUTdYLnD2wFktrj1uPpQSXs1fDyTBTz46+vl3V5zinZEpY5YN/K9Vx
1YJMxHcCjxC0KgPtxR6u2S2qUkwJcITThM/DTLwfp3KD8UXwuaELQXhIoxcE7sruz4rhNbQXKOHS
sUUMVPAszeIPC0cw21HY4yD/GVClrDHC06zJRUnZ7KuTeMruGtigVlSPb+Xk2vY5UoUHIQNQ2ytZ
sVdHKGr7h/ezs3ezrtsW516+7y6CIqtKBh2DHnF4Y+3u/8G699xn6p9seZTOkQJf8sAPPD9jvIlq
+pI3GjfN63H/YNS50R8nobd04IcwYG67R9J+x8zv1rQdz2aSVYOoflpeeik4onhixxNLBSNu4W+/
UnV8/OMsEh0Ar1MDaGXBHvRKw32jVUFu0pa4H8qij8WkSLx02c7CnHVRhuLSLkDVPVTTLFI23L+y
Ja6kkZnt+/HYQjtglJG1YkJOrNdOrLU29+P2S7MVwAq7Xe/mJ50OYXOQZ/PZ17HdCJF0EOM98LP5
D88RXRvmBA3HT14oGqLahEbBfF2yGzfi4TJ21XXGhULTHtSIalZog1JeFWDQxoT8q1PAAvyCVnc9
/hhAJJEp6+ZBCcjcl2EAOewMSWyfQHlkaVHuzloVl29e4gQyV6onLSr3UTLrK3rIvtJBKUKoP78k
bv/sczHHvfAXqUCr4ugWc6euR9cLeduyZprP8k5gb7KkHBsODvgziIAbP52VyDVQ6OVo48TSGApT
vmn45dh/EPrhMSKHs4najXcRe0sqtwxuPPqff4XI+ez8quxHY9Z/SKPlOgpr3lkpRHB+X8mPOQU4
V/xANuqzek0lk4pGS6GX5viW9thptGpQ1/l5EnexQgJUDpsPU2K6Qo8Ml57oM/eKuXomFCvzzx3o
jglyJ6N0x/XWbTJb4vWcSw8Et7/ERd7W91wV4VvDI3ktYzLjWhDtvxt2XLLYoIkvLyktdzgxwWFi
n0gpOCu5ANYAP+lIPtl3Lcg95Rwyy+GAq5LPnGRg5QtrpjfeaRFvkAW0RQJ3W65OvmmRcUwFrPOO
3lNkAROALxZ0oLg9w/VIR7PwUVbVp+ftvgT1oUiEiGEXCmBG0IewEFp6VDgjZLFG6auADlJsL93Z
GAO+5CuCFmQqAG/0+h0Kc8SWZSONrRPl7jubhhhW+0mrhDFb4AdM/RSNNSWH3+Qg7vN5hG3RugH5
9QjRK86CRaS5DkFMSnmtFGMpyrnPJNrI3gaUpmR7kYgBiUFEEDx6heIE/HIqXXtn+eVWKf0dk5kq
hLN2BAbZMZQBk2n+SVuzkM8LrBa1wCUL9vShl3GdRFL6ZkpDNqNI8CK7tuhVLUA/+L2kqXMHvozl
xGPewXOsNDQNQZxxN3wI6/FWJKLkEIUehjc0IAjvjbo5gqF1Pt/hL7kpLA/ifUKmpwaya3lLUIax
/QIWH3tOeBjfuJQOOe4keynNGVTg+OEom2FvtZ7KGvL5JCD1gw+qUz8j2SLZ2YJX2m8jBpwnGYDP
0z8QV9UfaCoGDaNucT4GpZDwUTTQx8I6SZJtdNTgONqtCg/C72D8UOtBp3TBv8ykUbCNEXkj/RBq
O3GKu3CExERO0QzPOJWpd8KHuN1ji9pu1S38Pz7gUAqhVcqsOZZFyIR2PSArpOY57YLpopI0aOBW
NRv3aCpNVbk5UBMWYFtdLEtlFX13frahrJQTuHrleXXXkt3HcpWyMMnFnshVgtv1u2+CBjICcjj3
WodYP73+ePhNh1nPkHIldj/wHDW3b63069XK3MT77kjaydqj2lQ/ebl39Ot43cPgcScQ4ZupBbJ8
KpirjInTNPhfpJTlrZYpTqU2HXIWJ7kJ92E5UvlwVzbA9CBrUxdezCfLITpdEPa9Zv6XRD6uHcjd
zS1meLnFqdatO9q5RFCDKLmaic1zKhK3oz4cSwbMSp5qC6JXR40LblEaFH8e+smbuCT8SdInCUns
d72Ltjcnk080rBdMSpq/7KUvE3x3vjWX/L2fsi78fVGu73hpsvb7/u8+X9Y9ny/A0PoTamdWZ2lo
ViwmR07c16ctEOaoKuzC+KxYNddXpUA+eyfQEYIVOLAP9V7Eh8T1M2yFne2Gir9er0eKjZjY8Xhl
SozTugycxUaI1n9390afIn6K51qnnCZeLYOX+qMvAwOM6j/dppQ8c0V+rzuAEZInX7j5+OXN++Au
pqDl6keDYKA9y5S40RA7EaUJ6/KSv4WHZ8CEoLmLfCHJqFO2bOABZL/K8533jinsmavvTcze/kH8
pqrjp2W39FpA7ql1OK2Yo8tPX2SVIlwo2jKlR0WgNZpMwiQm/0X+Pl7YV+SQaNoaqF+whNzZDjBL
4wEsdq65CG/APKotHrme+3nscqOMTyz5Z8vFOy3XTGuQhZ/RipGnwTS85LFPJbqEOAfyYR7wIuLO
Z2Fbb/hdegXO2QkFFZ7HrFsNXUtKWo83St06sJ4xpODUd8lh0zjEWp5OZ5tM5H4ZfBb/4F5uIQS1
Yz/q0vRG6KCKCTkqNmgEY5g4jKQgRblU1CzaMnlEXnI3e695d/lBshgovniE8Cw48ClJk2XbJjoD
uRDHS7x6nvDjtdQRwslXfhzwaP2Yg7EMXl/3LNXZ9v0G3VoXqIq+gq7VnoLaQ5/W0o56l0OLiqSt
XuF0RhtJ0rPp9nZBxebg/TcLzZNBs5RrXuVruP2jY0+d2kozgzkh0wBr8ifhLWHTe/3fOR1nfOpq
pfNyqgOUY0NIrxyr6UtTFPpkJh4YAF1nU+cmd2xh6Vl8t6DEeyW8jJOaM+7pYY7H73HAiGRACvxz
i1F9lQJMGAakGai/9jigPjWtHMvciTVBYjszFw+7FNGCPejI9Xu6UdU8xaOBTVwYhw9xyZum8+7n
qBgntW5+gSXs32KuTY9KhCpQtNnAwBbgnuksZTrqj0TEqTUc5yQRzMRoGc1bSOCQZe/5km8K3Ydq
xmaVokdo8Odr/mUlgMk8A8Vy/XdOBYzdUjXcYURR8tZnhYjLWj85dOjGF+Te1xNhCRRW+jdGUTEY
G3XfumOU31g+JfO6KXoNZAOZ66U262nnd++JA60+SYJbqmG17E8PEKLc4jXIb1l4zIesrwjBa5hV
68ManfGY3TIFqbs/uDkHYTv5AY+yvMEAmlNTJWiGzg+S1yR08kFsatrXfHXysEzDXju23sga0Lva
HnuWapMa0mnZgZ6d7NJwry3Bc0vM0Cj/yrEfijaiI8BxnRJPT8csNFum3cX1SdJmRJPabrnx+p5T
sq5/gCPR6n7Ax8+3VtDerU9Da3kAgHUC32220f1Jk7Vl4q5ggyOhHJIt0TAqgBu7Lbvuym4PGpfn
wtmRKDyMUb693svrQAw3jdgriT8XqgctyvfNhjG5lIH192XEXFcSXeFTU/IMeXe3jyPG1m9l3Hkg
QaCoKyPYyusTRZaTGMxmlhzO87nYnhQ3WkUouSMt4jwWYQCNcEgHLh0CT33/wnDf9d4ZGIGC17EF
fAwywMMic85o7gWYoH07h9Y1AbIZdraFrn8DTbPszYurG4QUqnaL0hOmsE0suvDrFB5uFNOx+dqt
YviPQW5QAIzh6P6ZwAYYMUOSh6dKRvmDNSFgjd5cVhcdPk36cJ4JX8w88N3QHTdq9vEcHTNwbeHo
5Fj0OL0tsZWmV+z6xog6hJSAvVSwWMkeweeuCZ9CDtnRkBNKVhOVPgnbx7Po1mVA49Bq6juHcln+
kW5csvWvuSqhUyhZcjWrj3rWRbqwCYN/oKSx0pVNNQGXCtiG+OE2B9RlmH1lgX3myJQM1u8SnEDV
prPARtKBJp/lIQtI2c4jwzPdBIW5I5AQXSbkzZVQO7z9OLuSINV/v67W8vUpcvgYMHT8fWxnI+hg
r0KbFk6NUEpkSvORyd5wgkeKpj/yM08xSIJKkblird1zZmz2HPqZmll8yMR2WCmU/03tYveZR5Kc
QRrOaJehC9TpHGqMAp+b//to5LqrvqRGDXL1pAkCTtFDBgxDW+7nyle0ybDZhCYN1Wzk8gc2aF4r
MljH0es8lsoBXnv+6kkv8MQ/Ef7vi9T/aKP3hhwfg9VZRQvpaUp4p3XxTcBwEbXR4OVVQScVxzce
IHhAw6xwwRwVnxITl6LQtqeUUHs2kph3BiQNP7VYTafQ1yvA/ULnmvgAdCk7N8UfE4PvevQGDHXz
pV4W/bqpAgsxr/XDthW/kQ32/iWsqyzTeP2dsRzdqrTmWE9T+taRt+u7614yWBYKsWGywruJ/Lbp
HQ3UeF1o66rMxo+gRBeFWsQqN/jjP6ehhsW3rgTL5x5WvAt2mwHYJ02tn5eCJjeDZ+Jp+Hy+TtVs
Ne+GFsVAQSV3USaD45573HZTLuAv0TzWWUfch7U+HrA9alQE83IBNcelTYBWi4Ca7yxm0u3hsL7a
q/+4EjPDm0sQB16+/n6UcocV6MRKLjrll2+hLagl3B+dxUMUMh55DFm7qUtcfq7bD7Irdp2cSOQg
S12RVJ2mWhiXNMpOQ8f1tzpBHSxlRAInn3riGKihwVJ+kfzNXNGDES0LXyawkEmuuu0Wo8IDE8eR
CSDGl1hcNCuk6GdvCCMf9Uk2w7Hm6GNPIclCArbWARagdbkwSwf9EgosMNBOlpzxZenz6j9yS4Fn
VdT/o0SsNdvmw28/9RUeEs4EoLBVRSxJ+7gU1k4nABZhpUWaGb1XG1FZcxgnRUL1msWkDcCMhmsz
7qIB/rYRkKLdLSn70dsjjWtgDh75cW2gyEOHA7hOExcqcRpfNCKwuzI2u4JiYG64fsU2eM2Yu+xs
gw8YIU2cR+DdivHTEIqjM/kk6W9IGullaKzlo1+Uaj5RGnx5oXEfs8wzyb2dm3e4Dyo0Q+Rv9PrC
kFG17T9CMFS9S00wtGLwrWqgASbxUCKhSzmP+opP6EB4EZtYFZksSzptM3s+qaItrQsZYu2XXeZU
4112QKMZdLZ7xG6uTusduasEGzHQ0e2vivLUzzfIJkyZ/ztZMUu/qa9EiS1TAuqAiXcXQgt8Z1SK
lMB7lOkpvXrt1ee2MxBuWWm2wPcwZsZtU+ZGRc1+BWs2A1R3gqlP5UIy9eaRG1ukWGwOy7+4khhi
PX1BKDtJsVnKWmkzIvupQq3pxwupExHXLV0jtq2xvpCujDWDqPz03gop4D6n6JxUZDvG2Jr5yt46
452h79El7eg/7xHFQ12wMMrsvs4+jticI3GQpHLVn3QFL9rRaQ9rYf02vFntsMtrVu5yRWKCMJbo
agSRPisWYdaMmLt4bF+cP6BAKO/bEETmv3ZaaY9EbwKbkPJdY9QFC7lZ2xy7ffBfBva9gD6/LRyP
JFA4oY/B68wAaEm0nJEThq8wtBmmaFwBuwoAtgzgbxs8Swg0f7Qbm1oamXWX8yObJwua4e/Gw8dz
HlyuowhBesRtAW0NO2lXSvRBHdt7mWu2ogzLO7gxaT/BD+/Sid6nQk86gJxdODhuVl3ufQZLjxmY
XQ4Yd58807wrc7XjMoiTTKujaURCAyDCNvqswzPyeDpqJi41PwCGkeyQfk6KB59CCUqP6JseJzUj
YNRdMRAK/DXvXEnJr1iwVFlFgRo2KshkasW7yZOzDmLjAzM6QnWoCm+oJC/k3Wj6wn5j5hPykz9w
nSlgqYabVhhyU7Tf3s8FKP3slLiM9kZsQ4k6mmmgeNgg7XVzzUEt/mWHA6BgqXyb6otGf10FmDFP
368/LO2+bEk/wTVtXzQ+7MLd21CwBG4p0jCzse+G2Du66rs7idBSxRbUdG7nOCjbg0H3u/l3JSQd
mW76SfGhsSNT9mNca6sYAPOM0clLinpAA8KhaZFtne+VbMwTK5WETfudAjo3dxJJ3Tn2Wfm10A9D
Zvm0WN+9aTvn1gZh6ZMTbDVhG5av0UHXx0VSRXNRQgyN3AnFy6jhcTpMDO7k+i/1AappETHXIDxF
akxsgY1nJNz7A/Jm+a068naWKyhIv4pLyl//nWDPgEiLcqQNLa4NxpqMKNaata/mA5jtVj97hyYb
CnD4FhKtoU123NZGcEc2i5ck+hppT/G92U8vZ1vpt0QoUZ3XvvHkp0Qxd2QTaj0Vaqxmue/Gpok9
rY+h7gBNdTmACmbycJs1/5ovMuTbMTeDvsownMitGrpfCAHJAai6drgUoj87e41psmcxirO25ZDi
DQO4BjmBAFenj9t1KSjEjQFEiebRgR3KYfHOxu/7R8flliYOy1ty0vJY7SITUV3XvjUwxnOTK/rk
NkOlO42I/c3ANIu/9uXsvjzJuqWHuesozVUgHFk34h46+LMJsQp8zYtzcsmhOx3vQNYhLZDmHyDu
Ms+orr5hP3lEBtBlxi4BB/1VTel9XUWG2GHhISDAfRhhbyx//eQwWej7OwW055wctmJvHBPG5cxs
cBtm4F5tT4SZ5Pla2Z3wBSTlEdAh1/Bk3DKFga060nYujlMae4yJx70VjwgeBlXu0qTvwUCWoLj9
q+4eZDygKVdlrF1voheHmYIII6RJYk0uT7Egej5ZPYo4eFkt60Dcfsh9OaIyRAB4QiYqAmemrhwS
cTFHMiOs+si1aeWVTUFx/HcdLR+ZOuTAfXK+BtVmi5slhpQeCwlfzhGf33GcgLOgPohF3fekssF4
8fHGwPH+e6lVp+LRyaceVvFmYNWGyQKu0+UCu5JmBBYYavg3qCt9Q8yIMU8qmDVYc+OwReWAvbIY
rLvvzkG4etbeMWTnvZGjolrEG/y0G/V+nY1y4HNiT3opRxhiiplXOUoCNVOoaMlJdNFa8lJdeSd4
x5UUTibI3IOF0NuJjG+aLWsTEn97DJDUsuncIjVgXuraydQvhZK9/x4NB1nkkKpjB+zu1WA7RTsj
VuIW69fPBC1g+2x7EEz5IbMUIchmFDH7bdpzpcuZcXhWPpR+LP1CDazB9zZnQ4VK1xpjRbiWJ+6D
NUgfmSiaRSCtJayU4HTTLoBs9peHPG/nLo1xXCm4hZyARpTwg7JnMqJXJMk08eCKyTH4kOEn4TId
yt2kzBE9tXgjRdSi9yLe08siby9ioeXVdOmCdRU6VYDJxZvq21+MHpTt3Q2zb2h+g+GTEEM3h/oI
lef3jqFJCOs6fBN8CrSEbcCV/thkZY75e+ixjyBkXt43Dlk7tlGgBoSXZjMIWbqF3RB2IFfvoGin
xuOv64hGMQQyY3AMHrkp5f1s0oOxWKhD3JccTV5Dnfw4n+Bs9gR/VH4KBpIUNBoJZytzeTYHWO5R
kJfyTLngZFQAmzdi61Gcv/jBzOVp0zvnFRjiyon4mrnV0/HLbqNzzdARL6Bk6y/B+MzSfLHzdvKx
8be4bfGVVUix8k7s1LhEiGDKDSU1vjan48WQZe6j5eZ0ahg3g7T/dQmqePWiGEZfARNcpLEpHvu3
0BgacV/475QLBwg52bE5ps7oEkDoQ5FtB8hljJJ03BFCzc/FUHlv8JtpaaG1xetJp7TZtqtC5JwT
2EMm5r9PaR/ii4k1tGlhRpL/KFQDUncz8P9OxsNTWkypcadCeO3tpfJMm37JeYttrRvOrCiwMtvm
KFcMOdq53iDWHf4eWg6dvly6cyD3VkvHrIeeteXkIHS0V2d3xC6iY3rsqq1riztmTkhG0Ho8oVAa
GPTp3a2bsJjIERznHbf8XE+7Wp4sc60KYoUCKH4fKVHpwHch+3E4Vl4EtbU4fxlIMvyri1mowtQv
cA1ZedNujf9ihh07ndS72zrlBRqLiJaS4Wo0Wn7d4LkF+kTKKa/0mc1EAtPPBGuxME5Ae4SbDkHj
3PA6mTS+xJvWyEQx2sVul0XslcYwvWJQWJxa17vsPlm9PWUZzrvMuz8uOLMhiTXJ1NLfzlSEWJQP
Lqgo6zxGaaQ4Aut2Bmj+BFnSakqlFKgaVaEkvPLBwtS+LqHivs+XmKQ51ia2vl9zCPNGVl4lAdML
dTgoXJRLQRb9FwMu8AaLWGU8AAccZlRCpBsfId8u4zXbdyqE3yf9uJMSo+ysiIORVYo5KGfWsu8I
etshhuEWMTcuAccjRbj/pX9C0KBbOmWVhVCAVRLQ/ggPTcVgqJdp6xNpZnpGJDEtrQVoZZmvqvay
FNk2/cPl/goQgdv1s81dd5PhK4/izZuYB1UYYuhv3vktHU60+LAZphnnyhU7BBszA3stSHUXqWSs
H9tI9CrsVbt9IPJxvyabaG3oJ+Lw73tiUWVcb2imbGYvfJ5iRjoUsaFDStDFbOwUZ9U2Wi18VRMS
OiUMlmNby9SiLzQDEBH11UKKBaZ33l4g+AzXXLkJNAxEJlRe32U1FPPy3Ojon3GlSSRdCs39/vXQ
tdxUCaGlvfdGaL5Az1Kni1wST+tAB5K9Kl5bO2KgNfG4qO3vVup26YKAvQ4ZSaqj8aRxGYNVXqX0
j9Cbj1vAsqLs8/RjaWfdzBhGiw/ktLvCHitPJPQnkxp59U8C6U1bpsVKpQfYo57zuxsH/BtGLIs5
7FRCxN1TRiI0NgZdU6tXiPsUZUyf56Iu7eIy7R1A5HItAYzWcYxurwW0EJXv3PxPMfYvpYhrKRgs
iVNls5HOnhZyC2cD6VsGSwVH/O9l4za2iZS/jEnZMGr31kBJLwIz9Wak1nbfVdDZMSiipJsdYrgY
S1YRorHOvf6vAVbeNDEzWXGk0PRabMcTmYQN0mFOjOFs7cVvRVnpTwEhQ/bYHz7E3q2L/SkZ0/Mv
kQJHP1J/Tmf0xOqBTEpFB2d9bD+QsQ53zqDiqHtkJWe21GLgLF7bHjFwE8P41KiUyxa96WwbVjLx
+TbYvHnVhSfA+830tw3xKw2SxQNx9mRDFaehgiYVt/2S96ApELjR6bsxXmU5Iq/P6nCZMAWuuKs+
878tsml05j/Hg96MlgLVhRbXhiLbvr5ruQiMpLtOoZsXu1ICgxzQRVeCi6m1Nkg/
`pragma protect end_protected
